magic
tech scmos
timestamp 1701903893
<< polysilicon >>
rect 5 71 7 83
rect 23 71 25 90
rect 41 71 43 83
rect 49 71 51 73
rect 57 71 59 83
rect 65 71 67 73
rect 86 71 88 113
rect 104 71 106 131
rect 122 71 124 83
rect 130 71 132 73
rect 138 71 140 83
rect 146 71 148 73
rect 168 71 170 91
rect 176 71 178 91
rect 192 71 194 73
rect 219 71 221 113
rect 227 71 229 131
rect 243 71 245 73
rect 265 71 267 94
rect 273 71 275 73
rect 314 71 316 73
rect 5 21 7 63
rect 23 21 25 63
rect 41 25 43 55
rect 49 25 51 55
rect 57 25 59 55
rect 65 25 67 55
rect 86 21 88 63
rect 104 21 106 63
rect 122 25 124 55
rect 130 25 132 55
rect 138 25 140 55
rect 146 25 148 55
rect 168 25 170 63
rect 176 25 178 63
rect 192 21 194 63
rect 219 25 221 63
rect 227 25 229 63
rect 243 21 245 63
rect 265 25 267 63
rect 273 25 275 63
rect 314 21 316 63
rect 5 15 7 17
rect 23 -22 25 17
rect 41 15 43 17
rect 49 -22 51 17
rect 57 15 59 17
rect 65 -22 67 17
rect 86 15 88 17
rect 104 -22 106 17
rect 122 15 124 17
rect 130 -22 132 17
rect 138 15 140 17
rect 146 -22 148 17
rect 168 15 170 17
rect 176 15 178 17
rect 192 15 194 17
rect 219 15 221 17
rect 227 15 229 17
rect 243 15 245 17
rect 265 15 267 17
rect 273 -8 275 17
rect 314 15 316 17
<< ndiffusion >>
rect -6 17 5 21
rect 7 17 8 21
rect 22 17 23 21
rect 25 17 26 21
rect 40 17 41 25
rect 43 17 49 25
rect 51 17 52 25
rect 56 17 57 25
rect 59 17 65 25
rect 67 17 68 25
rect 85 17 86 21
rect 88 17 89 21
rect 103 17 104 21
rect 106 17 107 21
rect 121 17 122 25
rect 124 17 130 25
rect 132 17 133 25
rect 137 17 138 25
rect 140 17 146 25
rect 148 17 149 25
rect 167 17 168 25
rect 170 17 176 25
rect 178 17 179 25
rect 191 17 192 21
rect 194 17 195 21
rect 218 17 219 25
rect 221 17 227 25
rect 229 17 230 25
rect 242 17 243 21
rect 245 17 246 21
rect 264 17 265 25
rect 267 17 268 25
rect 272 17 273 25
rect 275 17 276 25
rect 313 17 314 21
rect 316 17 317 21
<< pdiffusion >>
rect 4 63 5 71
rect 7 63 8 71
rect 22 63 23 71
rect 25 63 26 71
rect 40 55 41 71
rect 43 63 44 71
rect 48 63 49 71
rect 43 55 49 63
rect 51 55 52 71
rect 56 55 57 71
rect 59 63 65 71
rect 59 55 60 63
rect 64 55 65 63
rect 67 55 68 71
rect 85 63 86 71
rect 88 63 89 71
rect 103 63 104 71
rect 106 63 107 71
rect 121 55 122 71
rect 124 63 125 71
rect 129 63 130 71
rect 124 55 130 63
rect 132 55 133 71
rect 137 55 138 71
rect 140 63 146 71
rect 140 55 141 63
rect 145 55 146 63
rect 148 55 149 71
rect 167 63 168 71
rect 170 63 171 71
rect 175 63 176 71
rect 178 63 179 71
rect 191 63 192 71
rect 194 63 195 71
rect 218 63 219 71
rect 221 63 222 71
rect 226 63 227 71
rect 229 63 230 71
rect 242 63 243 71
rect 245 63 246 71
rect 264 63 265 71
rect 267 63 273 71
rect 275 63 276 71
rect 313 63 314 71
rect 316 63 317 71
<< metal1 >>
rect 108 131 227 135
rect 89 113 218 117
rect 4 106 171 110
rect 4 87 8 106
rect 22 94 26 97
rect 167 95 171 106
rect 175 95 179 98
rect 257 94 264 98
rect 8 83 40 87
rect 53 83 56 87
rect 92 83 121 87
rect 134 83 137 87
rect 0 79 321 80
rect 0 75 14 79
rect 18 75 97 79
rect 101 75 171 79
rect 175 75 188 79
rect 192 75 222 79
rect 226 75 239 79
rect 243 75 268 79
rect 272 75 310 79
rect 314 75 321 79
rect 0 74 321 75
rect 0 71 4 74
rect 18 71 22 74
rect 44 71 48 74
rect 81 71 85 74
rect 99 71 103 74
rect 125 71 129 74
rect 163 71 167 74
rect 179 71 183 74
rect 8 48 12 63
rect 26 48 30 63
rect 40 55 52 59
rect 56 67 68 71
rect 60 43 64 55
rect 89 48 93 63
rect 107 48 111 63
rect 121 55 133 59
rect 137 67 149 71
rect 187 71 191 74
rect 214 71 218 74
rect 230 71 234 74
rect 238 71 242 74
rect 260 71 264 74
rect 309 71 313 74
rect 141 43 145 55
rect 171 48 175 63
rect 195 48 199 63
rect 222 48 226 63
rect 246 48 250 63
rect 276 48 280 63
rect 171 44 188 48
rect 8 21 12 43
rect 26 21 30 43
rect 52 39 82 43
rect 52 25 56 39
rect 89 21 93 43
rect 107 21 111 43
rect 133 39 155 43
rect 133 25 137 39
rect 179 25 183 44
rect -10 14 -6 17
rect 18 14 22 17
rect 36 14 40 17
rect 68 14 72 17
rect 81 14 85 17
rect 99 14 103 17
rect 117 14 121 17
rect 149 14 153 17
rect 222 44 239 48
rect 195 21 199 43
rect 230 25 234 44
rect 268 44 310 48
rect 246 21 250 43
rect 268 25 272 44
rect 317 21 321 63
rect 163 14 167 17
rect 187 14 191 17
rect 214 14 218 17
rect 238 14 242 17
rect 260 14 264 17
rect 276 14 280 17
rect 309 14 313 17
rect -10 13 321 14
rect -10 9 -9 13
rect -5 9 82 13
rect 86 9 164 13
rect 168 9 188 13
rect 192 9 215 13
rect 219 9 239 13
rect 243 9 261 13
rect 265 9 310 13
rect 314 9 321 13
rect -10 8 321 9
rect 268 -12 272 -8
rect 26 -26 48 -22
rect 61 -26 64 -22
rect 107 -26 129 -22
rect 142 -26 145 -22
<< metal2 >>
rect 27 98 175 102
rect 48 80 52 83
rect 129 80 133 83
rect 252 80 256 94
rect 27 76 52 80
rect 108 76 133 80
rect 196 76 256 80
rect 27 48 31 76
rect 108 48 112 76
rect 196 48 200 76
rect 9 12 13 43
rect 90 12 94 43
rect 9 8 60 12
rect 90 8 141 12
rect 56 -22 60 8
rect 137 -22 141 8
rect 247 -8 251 43
rect 247 -12 263 -8
<< ntransistor >>
rect 5 17 7 21
rect 23 17 25 21
rect 41 17 43 25
rect 49 17 51 25
rect 57 17 59 25
rect 65 17 67 25
rect 86 17 88 21
rect 104 17 106 21
rect 122 17 124 25
rect 130 17 132 25
rect 138 17 140 25
rect 146 17 148 25
rect 168 17 170 25
rect 176 17 178 25
rect 192 17 194 21
rect 219 17 221 25
rect 227 17 229 25
rect 243 17 245 21
rect 265 17 267 25
rect 273 17 275 25
rect 314 17 316 21
<< ptransistor >>
rect 5 63 7 71
rect 23 63 25 71
rect 41 55 43 71
rect 49 55 51 71
rect 57 55 59 71
rect 65 55 67 71
rect 86 63 88 71
rect 104 63 106 71
rect 122 55 124 71
rect 130 55 132 71
rect 138 55 140 71
rect 146 55 148 71
rect 168 63 170 71
rect 176 63 178 71
rect 192 63 194 71
rect 219 63 221 71
rect 227 63 229 71
rect 243 63 245 71
rect 265 63 267 71
rect 273 63 275 71
rect 314 63 316 71
<< polycontact >>
rect 104 131 108 135
rect 227 131 231 135
rect 85 113 89 117
rect 22 90 26 94
rect 4 83 8 87
rect 40 83 44 87
rect 56 83 60 87
rect 88 83 92 87
rect 218 113 222 117
rect 167 91 171 95
rect 175 91 179 95
rect 121 83 125 87
rect 137 83 141 87
rect 264 94 268 98
rect 19 44 23 48
rect 82 39 86 43
rect 188 44 192 48
rect 239 44 243 48
rect 310 44 314 48
rect 272 -12 276 -8
rect 22 -26 26 -22
rect 48 -26 52 -22
rect 64 -26 68 -22
rect 103 -26 107 -22
rect 129 -26 133 -22
rect 145 -26 149 -22
<< ndcontact >>
rect -10 17 -6 21
rect 8 17 12 21
rect 18 17 22 21
rect 26 17 30 21
rect 36 17 40 25
rect 52 17 56 25
rect 68 17 72 25
rect 81 17 85 21
rect 89 17 93 21
rect 99 17 103 21
rect 107 17 111 21
rect 117 17 121 25
rect 133 17 137 25
rect 149 17 153 25
rect 163 17 167 25
rect 179 17 183 25
rect 187 17 191 21
rect 195 17 199 21
rect 214 17 218 25
rect 230 17 234 25
rect 238 17 242 21
rect 246 17 250 21
rect 260 17 264 25
rect 268 17 272 25
rect 276 17 280 25
rect 309 17 313 21
rect 317 17 321 21
<< pdcontact >>
rect 0 63 4 71
rect 8 63 12 71
rect 18 63 22 71
rect 26 63 30 71
rect 36 55 40 71
rect 44 63 48 71
rect 52 55 56 71
rect 60 55 64 63
rect 68 55 72 71
rect 81 63 85 71
rect 89 63 93 71
rect 99 63 103 71
rect 107 63 111 71
rect 117 55 121 71
rect 125 63 129 71
rect 133 55 137 71
rect 141 55 145 63
rect 149 55 153 71
rect 163 63 167 71
rect 171 63 175 71
rect 179 63 183 71
rect 187 63 191 71
rect 195 63 199 71
rect 214 63 218 71
rect 222 63 226 71
rect 230 63 234 71
rect 238 63 242 71
rect 246 63 250 71
rect 260 63 264 71
rect 276 63 280 71
rect 309 63 313 71
rect 317 63 321 71
<< m2contact >>
rect 22 97 27 102
rect 175 98 180 103
rect 252 94 257 99
rect 48 83 53 88
rect 129 83 134 88
rect 8 43 13 48
rect 26 43 31 48
rect 89 43 94 48
rect 107 43 112 48
rect 195 43 200 48
rect 246 43 251 48
rect 263 -13 268 -8
rect 56 -27 61 -22
rect 137 -27 142 -22
<< psubstratepcontact >>
rect -9 9 -5 13
rect 82 9 86 13
rect 164 9 168 13
rect 188 9 192 13
rect 215 9 219 13
rect 239 9 243 13
rect 261 9 265 13
rect 310 9 314 13
<< nsubstratencontact >>
rect 14 75 18 79
rect 97 75 101 79
rect 171 75 175 79
rect 188 75 192 79
rect 222 75 226 79
rect 239 75 243 79
rect 268 75 272 79
rect 310 75 314 79
<< labels >>
rlabel metal1 115 77 115 77 5 vdd
rlabel metal1 115 11 115 11 1 gnd
rlabel metal1 152 41 152 41 1 S
rlabel polycontact 6 85 6 85 1 A
rlabel polycontact 21 46 21 46 1 B
rlabel m2contact 10 45 10 45 1 not1_1
rlabel m2contact 28 45 28 45 1 not1_2
rlabel m2contact 91 46 91 46 1 not2_1
rlabel m2contact 109 45 109 45 1 not2_2
rlabel polycontact 84 41 84 41 1 out_XOR1
rlabel polycontact 190 46 190 46 1 out_AND1
rlabel polycontact 241 46 241 46 1 out_AND2
rlabel polycontact 106 133 106 133 5 cin
rlabel polycontact 312 46 312 46 1 out_OR
rlabel metal1 319 46 319 46 7 cout
<< end >>
