magic
tech scmos
timestamp 1701990606
<< polysilicon >>
rect -523 273 -521 275
rect -504 273 -502 275
rect -485 273 -483 303
rect -463 273 -461 275
rect -441 273 -439 275
rect -425 273 -423 294
rect -389 273 -387 294
rect -367 273 -365 275
rect -345 273 -343 275
rect -329 273 -327 303
rect -298 273 -296 275
rect -273 273 -271 275
rect -254 273 -252 303
rect -232 273 -230 275
rect -210 273 -208 275
rect -194 273 -192 294
rect -158 273 -156 294
rect -136 273 -134 275
rect -114 273 -112 275
rect -98 273 -96 303
rect -67 273 -65 275
rect 22 273 24 275
rect 41 273 43 303
rect 63 273 65 275
rect 85 273 87 275
rect 101 273 103 294
rect 137 273 139 294
rect 159 273 161 275
rect 181 273 183 275
rect 197 273 199 303
rect 228 273 230 275
rect 360 273 362 275
rect 379 273 381 303
rect 401 273 403 275
rect 423 273 425 275
rect 439 273 441 294
rect 475 273 477 294
rect 497 273 499 275
rect 519 273 521 275
rect 535 273 537 303
rect 566 273 568 275
rect 613 273 615 275
rect 632 273 634 303
rect 654 273 656 275
rect 676 273 678 275
rect 692 273 694 294
rect 728 273 730 294
rect 750 273 752 275
rect 772 273 774 275
rect 788 273 790 303
rect 819 273 821 275
rect 877 273 879 275
rect 896 273 898 303
rect 918 273 920 275
rect 940 273 942 275
rect 956 273 958 294
rect 992 273 994 294
rect 1014 273 1016 275
rect 1036 273 1038 275
rect 1052 273 1054 303
rect 1083 273 1085 275
rect 1161 273 1163 275
rect 1180 273 1182 303
rect 1202 273 1204 275
rect 1224 273 1226 275
rect 1240 273 1242 294
rect 1276 273 1278 294
rect 1298 273 1300 275
rect 1320 273 1322 275
rect 1336 273 1338 303
rect 1367 273 1369 275
rect 1413 273 1415 275
rect 1432 273 1434 303
rect 1454 273 1456 275
rect 1476 273 1478 275
rect 1492 273 1494 294
rect 1528 273 1530 294
rect 1550 273 1552 275
rect 1572 273 1574 275
rect 1588 273 1590 303
rect 1619 273 1621 275
rect 1672 273 1674 275
rect 1691 273 1693 303
rect 1713 273 1715 275
rect 1735 273 1737 275
rect 1751 273 1753 294
rect 1787 273 1789 294
rect 1809 273 1811 275
rect 1831 273 1833 275
rect 1847 273 1849 303
rect 1878 273 1880 275
rect -523 230 -521 265
rect -504 230 -502 265
rect -485 263 -483 265
rect -463 234 -461 257
rect -485 230 -483 232
rect -441 230 -439 265
rect -425 263 -423 265
rect -389 263 -387 265
rect -367 234 -365 257
rect -425 230 -423 232
rect -389 230 -387 232
rect -345 230 -343 265
rect -329 263 -327 265
rect -329 230 -327 232
rect -298 230 -296 265
rect -273 230 -271 265
rect -254 263 -252 265
rect -232 234 -230 257
rect -254 230 -252 232
rect -210 230 -208 265
rect -194 263 -192 265
rect -158 263 -156 265
rect -136 234 -134 257
rect -194 230 -192 232
rect -158 230 -156 232
rect -114 230 -112 265
rect -98 263 -96 265
rect -98 230 -96 232
rect -67 230 -65 265
rect 22 230 24 265
rect 41 263 43 265
rect 63 234 65 257
rect 41 230 43 232
rect 85 230 87 265
rect 101 263 103 265
rect 137 263 139 265
rect 159 234 161 257
rect 101 230 103 232
rect 137 230 139 232
rect 181 230 183 265
rect 197 263 199 265
rect 197 230 199 232
rect 228 230 230 265
rect 360 230 362 265
rect 379 263 381 265
rect 401 234 403 257
rect 379 230 381 232
rect 423 230 425 265
rect 439 263 441 265
rect 475 263 477 265
rect 497 234 499 257
rect 439 230 441 232
rect 475 230 477 232
rect 519 230 521 265
rect 535 263 537 265
rect 535 230 537 232
rect 566 230 568 265
rect 613 230 615 265
rect 632 263 634 265
rect 654 234 656 257
rect 632 230 634 232
rect 676 230 678 265
rect 692 263 694 265
rect 728 263 730 265
rect 750 234 752 257
rect 692 230 694 232
rect 728 230 730 232
rect 772 230 774 265
rect 788 263 790 265
rect 788 230 790 232
rect 819 230 821 265
rect 877 230 879 265
rect 896 263 898 265
rect 918 234 920 257
rect 896 230 898 232
rect 940 230 942 265
rect 956 263 958 265
rect 992 263 994 265
rect 1014 234 1016 257
rect 956 230 958 232
rect 992 230 994 232
rect 1036 230 1038 265
rect 1052 263 1054 265
rect 1052 230 1054 232
rect 1083 230 1085 265
rect 1161 230 1163 265
rect 1180 263 1182 265
rect 1202 234 1204 257
rect 1180 230 1182 232
rect 1224 230 1226 265
rect 1240 263 1242 265
rect 1276 263 1278 265
rect 1298 234 1300 257
rect 1240 230 1242 232
rect 1276 230 1278 232
rect 1320 230 1322 265
rect 1336 263 1338 265
rect 1336 230 1338 232
rect 1367 230 1369 265
rect 1413 230 1415 265
rect 1432 263 1434 265
rect 1454 234 1456 257
rect 1432 230 1434 232
rect 1476 230 1478 265
rect 1492 263 1494 265
rect 1528 263 1530 265
rect 1550 234 1552 257
rect 1492 230 1494 232
rect 1528 230 1530 232
rect 1572 230 1574 265
rect 1588 263 1590 265
rect 1588 230 1590 232
rect 1619 230 1621 265
rect 1672 230 1674 265
rect 1691 263 1693 265
rect 1713 234 1715 257
rect 1691 230 1693 232
rect 1735 230 1737 265
rect 1751 263 1753 265
rect 1787 263 1789 265
rect 1809 234 1811 257
rect 1751 230 1753 232
rect 1787 230 1789 232
rect 1831 230 1833 265
rect 1847 263 1849 265
rect 1847 230 1849 232
rect 1878 230 1880 265
rect -523 224 -521 226
rect -504 224 -502 226
rect -485 193 -483 226
rect -463 224 -461 226
rect -441 224 -439 226
rect -425 184 -423 226
rect -389 184 -387 226
rect -367 224 -365 226
rect -345 224 -343 226
rect -329 193 -327 226
rect -298 224 -296 226
rect -273 224 -271 226
rect -254 193 -252 226
rect -232 224 -230 226
rect -210 224 -208 226
rect -194 184 -192 226
rect -158 184 -156 226
rect -136 224 -134 226
rect -114 224 -112 226
rect -98 193 -96 226
rect -67 224 -65 226
rect 22 224 24 226
rect 41 193 43 226
rect 63 224 65 226
rect 85 224 87 226
rect 101 184 103 226
rect 137 184 139 226
rect 159 224 161 226
rect 181 224 183 226
rect 197 193 199 226
rect 228 224 230 226
rect 360 224 362 226
rect 379 193 381 226
rect 401 224 403 226
rect 423 224 425 226
rect 439 184 441 226
rect 475 184 477 226
rect 497 224 499 226
rect 519 224 521 226
rect 535 193 537 226
rect 566 224 568 226
rect 613 224 615 226
rect 632 193 634 226
rect 654 224 656 226
rect 676 224 678 226
rect 692 184 694 226
rect 728 184 730 226
rect 750 224 752 226
rect 772 224 774 226
rect 788 193 790 226
rect 819 224 821 226
rect 877 224 879 226
rect 896 193 898 226
rect 918 224 920 226
rect 940 224 942 226
rect 956 184 958 226
rect 992 184 994 226
rect 1014 224 1016 226
rect 1036 224 1038 226
rect 1052 193 1054 226
rect 1083 224 1085 226
rect 1161 224 1163 226
rect 1180 193 1182 226
rect 1202 224 1204 226
rect 1224 224 1226 226
rect 1240 184 1242 226
rect 1276 184 1278 226
rect 1298 224 1300 226
rect 1320 224 1322 226
rect 1336 193 1338 226
rect 1367 224 1369 226
rect 1413 224 1415 226
rect 1432 193 1434 226
rect 1454 224 1456 226
rect 1476 224 1478 226
rect 1492 184 1494 226
rect 1528 184 1530 226
rect 1550 224 1552 226
rect 1572 224 1574 226
rect 1588 193 1590 226
rect 1619 224 1621 226
rect 1672 224 1674 226
rect 1691 193 1693 226
rect 1713 224 1715 226
rect 1735 224 1737 226
rect 1751 184 1753 226
rect 1787 184 1789 226
rect 1809 224 1811 226
rect 1831 224 1833 226
rect 1847 193 1849 226
rect 1878 224 1880 226
rect 6 106 8 119
rect 22 106 24 126
rect 38 106 40 119
rect 46 106 48 108
rect 54 106 56 119
rect 62 106 64 108
rect 81 106 83 118
rect 89 106 91 118
rect 107 106 109 108
rect 135 106 137 119
rect 151 106 153 133
rect 167 106 169 119
rect 175 106 177 108
rect 183 106 185 119
rect 191 106 193 108
rect 210 106 212 118
rect 218 106 220 118
rect 236 106 238 108
rect 263 106 265 118
rect 271 106 273 118
rect 289 106 291 108
rect 321 106 323 119
rect 337 106 339 149
rect 353 106 355 119
rect 361 106 363 108
rect 369 106 371 119
rect 377 106 379 108
rect 396 106 398 118
rect 404 106 406 118
rect 422 106 424 108
rect 450 106 452 119
rect 466 106 468 135
rect 482 106 484 119
rect 490 106 492 108
rect 498 106 500 119
rect 506 106 508 108
rect 525 106 527 118
rect 533 106 535 118
rect 551 106 553 108
rect 578 106 580 118
rect 586 106 588 118
rect 604 106 606 108
rect 885 106 887 119
rect 901 106 903 145
rect 917 106 919 119
rect 925 106 927 108
rect 933 106 935 119
rect 941 106 943 108
rect 960 106 962 118
rect 968 106 970 118
rect 986 106 988 108
rect 1014 106 1016 119
rect 1030 106 1032 135
rect 1046 106 1048 119
rect 1054 106 1056 108
rect 1062 106 1064 119
rect 1070 106 1072 108
rect 1089 106 1091 118
rect 1097 106 1099 118
rect 1115 106 1117 108
rect 1142 106 1144 118
rect 1150 106 1152 118
rect 1168 106 1170 108
rect 1468 106 1470 119
rect 1484 106 1486 144
rect 1500 106 1502 119
rect 1508 106 1510 108
rect 1516 106 1518 119
rect 1524 106 1526 108
rect 1543 106 1545 118
rect 1551 106 1553 118
rect 1569 106 1571 108
rect 1597 106 1599 119
rect 1613 106 1615 135
rect 1629 106 1631 119
rect 1637 106 1639 108
rect 1645 106 1647 119
rect 1653 106 1655 108
rect 1672 106 1674 118
rect 1680 106 1682 118
rect 1698 106 1700 108
rect 1725 106 1727 118
rect 1733 106 1735 118
rect 1751 106 1753 108
rect 6 38 8 98
rect 22 38 24 98
rect 38 42 40 90
rect 46 42 48 90
rect 54 42 56 90
rect 62 42 64 90
rect 81 42 83 98
rect 89 42 91 98
rect 107 38 109 98
rect 135 38 137 98
rect 151 38 153 98
rect 167 42 169 90
rect 175 42 177 90
rect 183 42 185 90
rect 191 42 193 90
rect 210 42 212 98
rect 218 42 220 98
rect 236 38 238 98
rect 263 43 265 98
rect 271 43 273 98
rect 289 38 291 98
rect 321 38 323 98
rect 337 38 339 98
rect 353 42 355 90
rect 361 42 363 90
rect 369 42 371 90
rect 377 42 379 90
rect 396 42 398 98
rect 404 42 406 98
rect 6 32 8 34
rect 22 21 24 34
rect 38 32 40 34
rect 46 21 48 34
rect 54 32 56 34
rect 62 21 64 34
rect 81 32 83 34
rect 89 22 91 34
rect 107 32 109 34
rect 135 32 137 34
rect 151 21 153 34
rect 167 32 169 34
rect 175 21 177 34
rect 183 32 185 34
rect 191 21 193 34
rect 210 32 212 34
rect 218 22 220 34
rect 236 32 238 34
rect 263 32 265 35
rect 271 22 273 35
rect 422 38 424 98
rect 450 38 452 98
rect 466 38 468 98
rect 482 42 484 90
rect 490 42 492 90
rect 498 42 500 90
rect 506 42 508 90
rect 525 42 527 98
rect 533 42 535 98
rect 551 38 553 98
rect 578 43 580 98
rect 586 43 588 98
rect 604 38 606 98
rect 885 38 887 98
rect 901 38 903 98
rect 917 42 919 90
rect 925 42 927 90
rect 933 42 935 90
rect 941 42 943 90
rect 960 42 962 98
rect 968 42 970 98
rect 289 32 291 34
rect 321 32 323 34
rect 337 21 339 34
rect 353 32 355 34
rect 361 21 363 34
rect 369 32 371 34
rect 377 21 379 34
rect 396 32 398 34
rect 404 22 406 34
rect 422 32 424 34
rect 450 32 452 34
rect 466 21 468 34
rect 482 32 484 34
rect 490 21 492 34
rect 498 32 500 34
rect 506 21 508 34
rect 525 32 527 34
rect 533 22 535 34
rect 551 32 553 34
rect 578 32 580 35
rect 586 22 588 35
rect 986 38 988 98
rect 1014 38 1016 98
rect 1030 38 1032 98
rect 1046 42 1048 90
rect 1054 42 1056 90
rect 1062 42 1064 90
rect 1070 42 1072 90
rect 1089 42 1091 98
rect 1097 42 1099 98
rect 1115 38 1117 98
rect 1142 43 1144 98
rect 1150 43 1152 98
rect 1168 38 1170 98
rect 1468 38 1470 98
rect 1484 38 1486 98
rect 1500 42 1502 90
rect 1508 42 1510 90
rect 1516 42 1518 90
rect 1524 42 1526 90
rect 1543 42 1545 98
rect 1551 42 1553 98
rect 604 32 606 34
rect 885 32 887 34
rect 901 21 903 34
rect 917 32 919 34
rect 925 21 927 34
rect 933 32 935 34
rect 941 21 943 34
rect 960 32 962 34
rect 968 22 970 34
rect 986 32 988 34
rect 1014 32 1016 34
rect 1030 21 1032 34
rect 1046 32 1048 34
rect 1054 21 1056 34
rect 1062 32 1064 34
rect 1070 21 1072 34
rect 1089 32 1091 34
rect 1097 22 1099 34
rect 1115 32 1117 34
rect 1142 32 1144 35
rect 1150 22 1152 35
rect 1569 38 1571 98
rect 1597 38 1599 98
rect 1613 38 1615 98
rect 1629 42 1631 90
rect 1637 42 1639 90
rect 1645 42 1647 90
rect 1653 42 1655 90
rect 1672 42 1674 98
rect 1680 42 1682 98
rect 1698 38 1700 98
rect 1725 43 1727 98
rect 1733 43 1735 98
rect 1751 38 1753 98
rect 1168 32 1170 34
rect 1468 32 1470 34
rect 1484 21 1486 34
rect 1500 32 1502 34
rect 1508 21 1510 34
rect 1516 32 1518 34
rect 1524 21 1526 34
rect 1543 32 1545 34
rect 1551 22 1553 34
rect 1569 32 1571 34
rect 1597 32 1599 34
rect 1613 21 1615 34
rect 1629 32 1631 34
rect 1637 21 1639 34
rect 1645 32 1647 34
rect 1653 21 1655 34
rect 1672 32 1674 34
rect 1680 22 1682 34
rect 1698 32 1700 34
rect 1725 32 1727 35
rect 1733 22 1735 35
rect 1751 32 1753 34
rect 10 -100 12 -57
rect 29 -100 31 -70
rect 51 -100 53 -98
rect 73 -100 75 -98
rect 89 -100 91 -79
rect 125 -100 127 -79
rect 147 -100 149 -98
rect 169 -100 171 -98
rect 185 -100 187 -70
rect 216 -100 218 -98
rect 256 -100 258 -98
rect 275 -100 277 -70
rect 297 -100 299 -98
rect 319 -100 321 -98
rect 335 -100 337 -79
rect 371 -100 373 -79
rect 393 -100 395 -98
rect 415 -100 417 -98
rect 431 -100 433 -70
rect 462 -100 464 -98
rect 757 -100 759 -98
rect 776 -100 778 -70
rect 798 -100 800 -98
rect 820 -100 822 -98
rect 836 -100 838 -79
rect 872 -100 874 -79
rect 894 -100 896 -98
rect 916 -100 918 -98
rect 932 -100 934 -70
rect 963 -100 965 -98
rect 1069 -100 1071 -98
rect 1088 -100 1090 -70
rect 1110 -100 1112 -98
rect 1132 -100 1134 -98
rect 1148 -100 1150 -79
rect 1184 -100 1186 -79
rect 1206 -100 1208 -98
rect 1228 -100 1230 -98
rect 1244 -100 1246 -70
rect 1275 -100 1277 -98
rect 1368 -100 1370 -98
rect 1387 -100 1389 -70
rect 1409 -100 1411 -98
rect 1431 -100 1433 -98
rect 1447 -100 1449 -79
rect 1483 -100 1485 -79
rect 1505 -100 1507 -98
rect 1527 -100 1529 -98
rect 1543 -100 1545 -70
rect 1574 -100 1576 -98
rect 10 -143 12 -108
rect 29 -110 31 -108
rect 51 -139 53 -116
rect 29 -143 31 -141
rect 73 -143 75 -108
rect 89 -110 91 -108
rect 125 -110 127 -108
rect 147 -139 149 -116
rect 89 -143 91 -141
rect 125 -143 127 -141
rect 169 -143 171 -108
rect 185 -110 187 -108
rect 185 -143 187 -141
rect 216 -143 218 -108
rect 256 -143 258 -108
rect 275 -110 277 -108
rect 297 -139 299 -116
rect 275 -143 277 -141
rect 319 -143 321 -108
rect 335 -110 337 -108
rect 371 -110 373 -108
rect 393 -139 395 -116
rect 335 -143 337 -141
rect 371 -143 373 -141
rect 415 -143 417 -108
rect 431 -110 433 -108
rect 431 -143 433 -141
rect 462 -143 464 -108
rect 757 -143 759 -108
rect 776 -110 778 -108
rect 798 -139 800 -116
rect 776 -143 778 -141
rect 820 -143 822 -108
rect 836 -110 838 -108
rect 872 -110 874 -108
rect 894 -139 896 -116
rect 836 -143 838 -141
rect 872 -143 874 -141
rect 916 -143 918 -108
rect 932 -110 934 -108
rect 932 -143 934 -141
rect 963 -143 965 -108
rect 1069 -143 1071 -108
rect 1088 -110 1090 -108
rect 1110 -139 1112 -116
rect 1088 -143 1090 -141
rect 1132 -143 1134 -108
rect 1148 -110 1150 -108
rect 1184 -110 1186 -108
rect 1206 -139 1208 -116
rect 1148 -143 1150 -141
rect 1184 -143 1186 -141
rect 1228 -143 1230 -108
rect 1244 -110 1246 -108
rect 1244 -143 1246 -141
rect 1275 -143 1277 -108
rect 1368 -143 1370 -108
rect 1387 -110 1389 -108
rect 1409 -139 1411 -116
rect 1387 -143 1389 -141
rect 1431 -143 1433 -108
rect 1447 -110 1449 -108
rect 1483 -110 1485 -108
rect 1505 -139 1507 -116
rect 1447 -143 1449 -141
rect 1483 -143 1485 -141
rect 1527 -143 1529 -108
rect 1543 -110 1545 -108
rect 1543 -143 1545 -141
rect 1574 -143 1576 -108
rect 10 -149 12 -147
rect 29 -180 31 -147
rect 51 -149 53 -147
rect 73 -149 75 -147
rect 89 -189 91 -147
rect 125 -189 127 -147
rect 147 -149 149 -147
rect 169 -149 171 -147
rect 185 -180 187 -147
rect 216 -149 218 -147
rect 256 -149 258 -147
rect 275 -180 277 -147
rect 297 -149 299 -147
rect 319 -149 321 -147
rect 335 -189 337 -147
rect 371 -189 373 -147
rect 393 -149 395 -147
rect 415 -149 417 -147
rect 431 -180 433 -147
rect 462 -149 464 -147
rect 757 -149 759 -147
rect 776 -180 778 -147
rect 798 -149 800 -147
rect 820 -149 822 -147
rect 836 -189 838 -147
rect 872 -189 874 -147
rect 894 -149 896 -147
rect 916 -149 918 -147
rect 932 -180 934 -147
rect 963 -149 965 -147
rect 1069 -149 1071 -147
rect 1088 -180 1090 -147
rect 1110 -149 1112 -147
rect 1132 -149 1134 -147
rect 1148 -189 1150 -147
rect 1184 -189 1186 -147
rect 1206 -149 1208 -147
rect 1228 -149 1230 -147
rect 1244 -180 1246 -147
rect 1275 -149 1277 -147
rect 1368 -149 1370 -147
rect 1387 -180 1389 -147
rect 1409 -149 1411 -147
rect 1431 -149 1433 -147
rect 1447 -189 1449 -147
rect 1483 -189 1485 -147
rect 1505 -149 1507 -147
rect 1527 -149 1529 -147
rect 1543 -180 1545 -147
rect 1574 -149 1576 -147
<< ndiffusion >>
rect -524 226 -523 230
rect -521 226 -520 230
rect -505 226 -504 230
rect -502 226 -501 230
rect -486 226 -485 230
rect -483 226 -482 230
rect -464 226 -463 234
rect -461 226 -460 234
rect -442 226 -441 230
rect -439 226 -438 230
rect -426 226 -425 230
rect -423 226 -422 230
rect -390 226 -389 230
rect -387 226 -386 230
rect -368 226 -367 234
rect -365 226 -364 234
rect -346 226 -345 230
rect -343 226 -342 230
rect -330 226 -329 230
rect -327 226 -326 230
rect -299 226 -298 230
rect -296 226 -295 230
rect -274 226 -273 230
rect -271 226 -270 230
rect -255 226 -254 230
rect -252 226 -251 230
rect -233 226 -232 234
rect -230 226 -229 234
rect -211 226 -210 230
rect -208 226 -207 230
rect -195 226 -194 230
rect -192 226 -191 230
rect -159 226 -158 230
rect -156 226 -155 230
rect -137 226 -136 234
rect -134 226 -133 234
rect -115 226 -114 230
rect -112 226 -111 230
rect -99 226 -98 230
rect -96 226 -95 230
rect -68 226 -67 230
rect -65 226 -64 230
rect 21 226 22 230
rect 24 226 25 230
rect 40 226 41 230
rect 43 226 44 230
rect 62 226 63 234
rect 65 226 66 234
rect 84 226 85 230
rect 87 226 88 230
rect 100 226 101 230
rect 103 226 104 230
rect 136 226 137 230
rect 139 226 140 230
rect 158 226 159 234
rect 161 226 162 234
rect 180 226 181 230
rect 183 226 184 230
rect 196 226 197 230
rect 199 226 200 230
rect 227 226 228 230
rect 230 226 231 230
rect 359 226 360 230
rect 362 226 363 230
rect 378 226 379 230
rect 381 226 382 230
rect 400 226 401 234
rect 403 226 404 234
rect 422 226 423 230
rect 425 226 426 230
rect 438 226 439 230
rect 441 226 442 230
rect 474 226 475 230
rect 477 226 478 230
rect 496 226 497 234
rect 499 226 500 234
rect 518 226 519 230
rect 521 226 522 230
rect 534 226 535 230
rect 537 226 538 230
rect 565 226 566 230
rect 568 226 569 230
rect 612 226 613 230
rect 615 226 616 230
rect 631 226 632 230
rect 634 226 635 230
rect 653 226 654 234
rect 656 226 657 234
rect 675 226 676 230
rect 678 226 679 230
rect 691 226 692 230
rect 694 226 695 230
rect 727 226 728 230
rect 730 226 731 230
rect 749 226 750 234
rect 752 226 753 234
rect 771 226 772 230
rect 774 226 775 230
rect 787 226 788 230
rect 790 226 791 230
rect 818 226 819 230
rect 821 226 822 230
rect 876 226 877 230
rect 879 226 880 230
rect 895 226 896 230
rect 898 226 899 230
rect 917 226 918 234
rect 920 226 921 234
rect 939 226 940 230
rect 942 226 943 230
rect 955 226 956 230
rect 958 226 959 230
rect 991 226 992 230
rect 994 226 995 230
rect 1013 226 1014 234
rect 1016 226 1017 234
rect 1035 226 1036 230
rect 1038 226 1039 230
rect 1051 226 1052 230
rect 1054 226 1055 230
rect 1082 226 1083 230
rect 1085 226 1086 230
rect 1160 226 1161 230
rect 1163 226 1164 230
rect 1179 226 1180 230
rect 1182 226 1183 230
rect 1201 226 1202 234
rect 1204 226 1205 234
rect 1223 226 1224 230
rect 1226 226 1227 230
rect 1239 226 1240 230
rect 1242 226 1243 230
rect 1275 226 1276 230
rect 1278 226 1279 230
rect 1297 226 1298 234
rect 1300 226 1301 234
rect 1319 226 1320 230
rect 1322 226 1323 230
rect 1335 226 1336 230
rect 1338 226 1339 230
rect 1366 226 1367 230
rect 1369 226 1370 230
rect 1412 226 1413 230
rect 1415 226 1416 230
rect 1431 226 1432 230
rect 1434 226 1435 230
rect 1453 226 1454 234
rect 1456 226 1457 234
rect 1475 226 1476 230
rect 1478 226 1479 230
rect 1491 226 1492 230
rect 1494 226 1495 230
rect 1527 226 1528 230
rect 1530 226 1531 230
rect 1549 226 1550 234
rect 1552 226 1553 234
rect 1571 226 1572 230
rect 1574 226 1575 230
rect 1587 226 1588 230
rect 1590 226 1591 230
rect 1618 226 1619 230
rect 1621 226 1622 230
rect 1671 226 1672 230
rect 1674 226 1675 230
rect 1690 226 1691 230
rect 1693 226 1694 230
rect 1712 226 1713 234
rect 1715 226 1716 234
rect 1734 226 1735 230
rect 1737 226 1738 230
rect 1750 226 1751 230
rect 1753 226 1754 230
rect 1786 226 1787 230
rect 1789 226 1790 230
rect 1808 226 1809 234
rect 1811 226 1812 234
rect 1830 226 1831 230
rect 1833 226 1834 230
rect 1846 226 1847 230
rect 1849 226 1850 230
rect 1877 226 1878 230
rect 1880 226 1881 230
rect 5 34 6 38
rect 8 34 9 38
rect 21 34 22 38
rect 24 34 25 38
rect 37 34 38 42
rect 40 34 46 42
rect 48 34 49 42
rect 53 34 54 42
rect 56 34 62 42
rect 64 34 65 42
rect 78 34 81 42
rect 83 34 89 42
rect 91 34 94 42
rect 106 34 107 38
rect 109 34 110 38
rect 134 34 135 38
rect 137 34 138 38
rect 150 34 151 38
rect 153 34 154 38
rect 166 34 167 42
rect 169 34 175 42
rect 177 34 178 42
rect 182 34 183 42
rect 185 34 191 42
rect 193 34 194 42
rect 207 34 210 42
rect 212 34 218 42
rect 220 34 223 42
rect 235 34 236 38
rect 238 34 239 38
rect 261 35 263 43
rect 265 35 266 43
rect 270 35 271 43
rect 273 35 274 43
rect 287 34 289 38
rect 291 34 293 38
rect 320 34 321 38
rect 323 34 324 38
rect 336 34 337 38
rect 339 34 340 38
rect 352 34 353 42
rect 355 34 361 42
rect 363 34 364 42
rect 368 34 369 42
rect 371 34 377 42
rect 379 34 380 42
rect 393 34 396 42
rect 398 34 404 42
rect 406 34 409 42
rect 421 34 422 38
rect 424 34 425 38
rect 449 34 450 38
rect 452 34 453 38
rect 465 34 466 38
rect 468 34 469 38
rect 481 34 482 42
rect 484 34 490 42
rect 492 34 493 42
rect 497 34 498 42
rect 500 34 506 42
rect 508 34 509 42
rect 522 34 525 42
rect 527 34 533 42
rect 535 34 538 42
rect 550 34 551 38
rect 553 34 554 38
rect 576 35 578 43
rect 580 35 581 43
rect 585 35 586 43
rect 588 35 589 43
rect 602 34 604 38
rect 606 34 608 38
rect 884 34 885 38
rect 887 34 888 38
rect 900 34 901 38
rect 903 34 904 38
rect 916 34 917 42
rect 919 34 925 42
rect 927 34 928 42
rect 932 34 933 42
rect 935 34 941 42
rect 943 34 944 42
rect 957 34 960 42
rect 962 34 968 42
rect 970 34 973 42
rect 985 34 986 38
rect 988 34 989 38
rect 1013 34 1014 38
rect 1016 34 1017 38
rect 1029 34 1030 38
rect 1032 34 1033 38
rect 1045 34 1046 42
rect 1048 34 1054 42
rect 1056 34 1057 42
rect 1061 34 1062 42
rect 1064 34 1070 42
rect 1072 34 1073 42
rect 1086 34 1089 42
rect 1091 34 1097 42
rect 1099 34 1102 42
rect 1114 34 1115 38
rect 1117 34 1118 38
rect 1140 35 1142 43
rect 1144 35 1145 43
rect 1149 35 1150 43
rect 1152 35 1153 43
rect 1166 34 1168 38
rect 1170 34 1172 38
rect 1467 34 1468 38
rect 1470 34 1471 38
rect 1483 34 1484 38
rect 1486 34 1487 38
rect 1499 34 1500 42
rect 1502 34 1508 42
rect 1510 34 1511 42
rect 1515 34 1516 42
rect 1518 34 1524 42
rect 1526 34 1527 42
rect 1540 34 1543 42
rect 1545 34 1551 42
rect 1553 34 1556 42
rect 1568 34 1569 38
rect 1571 34 1572 38
rect 1596 34 1597 38
rect 1599 34 1600 38
rect 1612 34 1613 38
rect 1615 34 1616 38
rect 1628 34 1629 42
rect 1631 34 1637 42
rect 1639 34 1640 42
rect 1644 34 1645 42
rect 1647 34 1653 42
rect 1655 34 1656 42
rect 1669 34 1672 42
rect 1674 34 1680 42
rect 1682 34 1685 42
rect 1697 34 1698 38
rect 1700 34 1701 38
rect 1723 35 1725 43
rect 1727 35 1728 43
rect 1732 35 1733 43
rect 1735 35 1736 43
rect 1749 34 1751 38
rect 1753 34 1755 38
rect 9 -147 10 -143
rect 12 -147 13 -143
rect 28 -147 29 -143
rect 31 -147 32 -143
rect 50 -147 51 -139
rect 53 -147 54 -139
rect 72 -147 73 -143
rect 75 -147 76 -143
rect 88 -147 89 -143
rect 91 -147 92 -143
rect 124 -147 125 -143
rect 127 -147 128 -143
rect 146 -147 147 -139
rect 149 -147 150 -139
rect 168 -147 169 -143
rect 171 -147 172 -143
rect 184 -147 185 -143
rect 187 -147 188 -143
rect 215 -147 216 -143
rect 218 -147 219 -143
rect 255 -147 256 -143
rect 258 -147 259 -143
rect 274 -147 275 -143
rect 277 -147 278 -143
rect 296 -147 297 -139
rect 299 -147 300 -139
rect 318 -147 319 -143
rect 321 -147 322 -143
rect 334 -147 335 -143
rect 337 -147 338 -143
rect 370 -147 371 -143
rect 373 -147 374 -143
rect 392 -147 393 -139
rect 395 -147 396 -139
rect 414 -147 415 -143
rect 417 -147 418 -143
rect 430 -147 431 -143
rect 433 -147 434 -143
rect 461 -147 462 -143
rect 464 -147 465 -143
rect 756 -147 757 -143
rect 759 -147 760 -143
rect 775 -147 776 -143
rect 778 -147 779 -143
rect 797 -147 798 -139
rect 800 -147 801 -139
rect 819 -147 820 -143
rect 822 -147 823 -143
rect 835 -147 836 -143
rect 838 -147 839 -143
rect 871 -147 872 -143
rect 874 -147 875 -143
rect 893 -147 894 -139
rect 896 -147 897 -139
rect 915 -147 916 -143
rect 918 -147 919 -143
rect 931 -147 932 -143
rect 934 -147 935 -143
rect 962 -147 963 -143
rect 965 -147 966 -143
rect 1068 -147 1069 -143
rect 1071 -147 1072 -143
rect 1087 -147 1088 -143
rect 1090 -147 1091 -143
rect 1109 -147 1110 -139
rect 1112 -147 1113 -139
rect 1131 -147 1132 -143
rect 1134 -147 1135 -143
rect 1147 -147 1148 -143
rect 1150 -147 1151 -143
rect 1183 -147 1184 -143
rect 1186 -147 1187 -143
rect 1205 -147 1206 -139
rect 1208 -147 1209 -139
rect 1227 -147 1228 -143
rect 1230 -147 1231 -143
rect 1243 -147 1244 -143
rect 1246 -147 1247 -143
rect 1274 -147 1275 -143
rect 1277 -147 1278 -143
rect 1367 -147 1368 -143
rect 1370 -147 1371 -143
rect 1386 -147 1387 -143
rect 1389 -147 1390 -143
rect 1408 -147 1409 -139
rect 1411 -147 1412 -139
rect 1430 -147 1431 -143
rect 1433 -147 1434 -143
rect 1446 -147 1447 -143
rect 1449 -147 1450 -143
rect 1482 -147 1483 -143
rect 1485 -147 1486 -143
rect 1504 -147 1505 -139
rect 1507 -147 1508 -139
rect 1526 -147 1527 -143
rect 1529 -147 1530 -143
rect 1542 -147 1543 -143
rect 1545 -147 1546 -143
rect 1573 -147 1574 -143
rect 1576 -147 1577 -143
<< pdiffusion >>
rect -524 265 -523 273
rect -521 265 -520 273
rect -505 265 -504 273
rect -502 265 -501 273
rect -486 265 -485 273
rect -483 265 -482 273
rect -464 257 -463 273
rect -461 257 -460 273
rect -442 265 -441 273
rect -439 265 -438 273
rect -426 265 -425 273
rect -423 265 -422 273
rect -390 265 -389 273
rect -387 265 -386 273
rect -368 257 -367 273
rect -365 257 -364 273
rect -346 265 -345 273
rect -343 265 -342 273
rect -330 265 -329 273
rect -327 265 -326 273
rect -299 265 -298 273
rect -296 265 -295 273
rect -274 265 -273 273
rect -271 265 -270 273
rect -255 265 -254 273
rect -252 265 -251 273
rect -233 257 -232 273
rect -230 257 -229 273
rect -211 265 -210 273
rect -208 265 -207 273
rect -195 265 -194 273
rect -192 265 -191 273
rect -159 265 -158 273
rect -156 265 -155 273
rect -137 257 -136 273
rect -134 257 -133 273
rect -115 265 -114 273
rect -112 265 -111 273
rect -99 265 -98 273
rect -96 265 -95 273
rect -68 265 -67 273
rect -65 265 -64 273
rect 21 265 22 273
rect 24 265 25 273
rect 40 265 41 273
rect 43 265 44 273
rect 62 257 63 273
rect 65 257 66 273
rect 84 265 85 273
rect 87 265 88 273
rect 100 265 101 273
rect 103 265 104 273
rect 136 265 137 273
rect 139 265 140 273
rect 158 257 159 273
rect 161 257 162 273
rect 180 265 181 273
rect 183 265 184 273
rect 196 265 197 273
rect 199 265 200 273
rect 227 265 228 273
rect 230 265 231 273
rect 359 265 360 273
rect 362 265 363 273
rect 378 265 379 273
rect 381 265 382 273
rect 400 257 401 273
rect 403 257 404 273
rect 422 265 423 273
rect 425 265 426 273
rect 438 265 439 273
rect 441 265 442 273
rect 474 265 475 273
rect 477 265 478 273
rect 496 257 497 273
rect 499 257 500 273
rect 518 265 519 273
rect 521 265 522 273
rect 534 265 535 273
rect 537 265 538 273
rect 565 265 566 273
rect 568 265 569 273
rect 612 265 613 273
rect 615 265 616 273
rect 631 265 632 273
rect 634 265 635 273
rect 653 257 654 273
rect 656 257 657 273
rect 675 265 676 273
rect 678 265 679 273
rect 691 265 692 273
rect 694 265 695 273
rect 727 265 728 273
rect 730 265 731 273
rect 749 257 750 273
rect 752 257 753 273
rect 771 265 772 273
rect 774 265 775 273
rect 787 265 788 273
rect 790 265 791 273
rect 818 265 819 273
rect 821 265 822 273
rect 876 265 877 273
rect 879 265 880 273
rect 895 265 896 273
rect 898 265 899 273
rect 917 257 918 273
rect 920 257 921 273
rect 939 265 940 273
rect 942 265 943 273
rect 955 265 956 273
rect 958 265 959 273
rect 991 265 992 273
rect 994 265 995 273
rect 1013 257 1014 273
rect 1016 257 1017 273
rect 1035 265 1036 273
rect 1038 265 1039 273
rect 1051 265 1052 273
rect 1054 265 1055 273
rect 1082 265 1083 273
rect 1085 265 1086 273
rect 1160 265 1161 273
rect 1163 265 1164 273
rect 1179 265 1180 273
rect 1182 265 1183 273
rect 1201 257 1202 273
rect 1204 257 1205 273
rect 1223 265 1224 273
rect 1226 265 1227 273
rect 1239 265 1240 273
rect 1242 265 1243 273
rect 1275 265 1276 273
rect 1278 265 1279 273
rect 1297 257 1298 273
rect 1300 257 1301 273
rect 1319 265 1320 273
rect 1322 265 1323 273
rect 1335 265 1336 273
rect 1338 265 1339 273
rect 1366 265 1367 273
rect 1369 265 1370 273
rect 1412 265 1413 273
rect 1415 265 1416 273
rect 1431 265 1432 273
rect 1434 265 1435 273
rect 1453 257 1454 273
rect 1456 257 1457 273
rect 1475 265 1476 273
rect 1478 265 1479 273
rect 1491 265 1492 273
rect 1494 265 1495 273
rect 1527 265 1528 273
rect 1530 265 1531 273
rect 1549 257 1550 273
rect 1552 257 1553 273
rect 1571 265 1572 273
rect 1574 265 1575 273
rect 1587 265 1588 273
rect 1590 265 1591 273
rect 1618 265 1619 273
rect 1621 265 1622 273
rect 1671 265 1672 273
rect 1674 265 1675 273
rect 1690 265 1691 273
rect 1693 265 1694 273
rect 1712 257 1713 273
rect 1715 257 1716 273
rect 1734 265 1735 273
rect 1737 265 1738 273
rect 1750 265 1751 273
rect 1753 265 1754 273
rect 1786 265 1787 273
rect 1789 265 1790 273
rect 1808 257 1809 273
rect 1811 257 1812 273
rect 1830 265 1831 273
rect 1833 265 1834 273
rect 1846 265 1847 273
rect 1849 265 1850 273
rect 1877 265 1878 273
rect 1880 265 1881 273
rect 5 98 6 106
rect 8 98 9 106
rect 21 98 22 106
rect 24 98 25 106
rect 37 90 38 106
rect 40 98 41 106
rect 45 98 46 106
rect 40 90 46 98
rect 48 90 49 106
rect 53 90 54 106
rect 56 98 62 106
rect 56 90 57 98
rect 61 90 62 98
rect 64 90 65 106
rect 74 104 81 106
rect 74 100 75 104
rect 79 100 81 104
rect 74 98 81 100
rect 83 104 89 106
rect 83 100 84 104
rect 88 100 89 104
rect 83 98 89 100
rect 91 104 98 106
rect 91 100 93 104
rect 97 100 98 104
rect 91 98 98 100
rect 106 98 107 106
rect 109 98 110 106
rect 134 98 135 106
rect 137 98 138 106
rect 150 98 151 106
rect 153 98 154 106
rect 166 90 167 106
rect 169 98 170 106
rect 174 98 175 106
rect 169 90 175 98
rect 177 90 178 106
rect 182 90 183 106
rect 185 98 191 106
rect 185 90 186 98
rect 190 90 191 98
rect 193 90 194 106
rect 203 104 210 106
rect 203 100 204 104
rect 208 100 210 104
rect 203 98 210 100
rect 212 104 218 106
rect 212 100 213 104
rect 217 100 218 104
rect 212 98 218 100
rect 220 104 227 106
rect 220 100 222 104
rect 226 100 227 104
rect 220 98 227 100
rect 235 98 236 106
rect 238 98 239 106
rect 261 98 263 106
rect 265 98 271 106
rect 273 98 274 106
rect 287 98 289 106
rect 291 98 293 106
rect 320 98 321 106
rect 323 98 324 106
rect 336 98 337 106
rect 339 98 340 106
rect 352 90 353 106
rect 355 98 356 106
rect 360 98 361 106
rect 355 90 361 98
rect 363 90 364 106
rect 368 90 369 106
rect 371 98 377 106
rect 371 90 372 98
rect 376 90 377 98
rect 379 90 380 106
rect 389 104 396 106
rect 389 100 390 104
rect 394 100 396 104
rect 389 98 396 100
rect 398 104 404 106
rect 398 100 399 104
rect 403 100 404 104
rect 398 98 404 100
rect 406 104 413 106
rect 406 100 408 104
rect 412 100 413 104
rect 406 98 413 100
rect 421 98 422 106
rect 424 98 425 106
rect 449 98 450 106
rect 452 98 453 106
rect 465 98 466 106
rect 468 98 469 106
rect 481 90 482 106
rect 484 98 485 106
rect 489 98 490 106
rect 484 90 490 98
rect 492 90 493 106
rect 497 90 498 106
rect 500 98 506 106
rect 500 90 501 98
rect 505 90 506 98
rect 508 90 509 106
rect 518 104 525 106
rect 518 100 519 104
rect 523 100 525 104
rect 518 98 525 100
rect 527 104 533 106
rect 527 100 528 104
rect 532 100 533 104
rect 527 98 533 100
rect 535 104 542 106
rect 535 100 537 104
rect 541 100 542 104
rect 535 98 542 100
rect 550 98 551 106
rect 553 98 554 106
rect 576 98 578 106
rect 580 98 586 106
rect 588 98 589 106
rect 602 98 604 106
rect 606 98 608 106
rect 884 98 885 106
rect 887 98 888 106
rect 900 98 901 106
rect 903 98 904 106
rect 916 90 917 106
rect 919 98 920 106
rect 924 98 925 106
rect 919 90 925 98
rect 927 90 928 106
rect 932 90 933 106
rect 935 98 941 106
rect 935 90 936 98
rect 940 90 941 98
rect 943 90 944 106
rect 953 104 960 106
rect 953 100 954 104
rect 958 100 960 104
rect 953 98 960 100
rect 962 104 968 106
rect 962 100 963 104
rect 967 100 968 104
rect 962 98 968 100
rect 970 104 977 106
rect 970 100 972 104
rect 976 100 977 104
rect 970 98 977 100
rect 985 98 986 106
rect 988 98 989 106
rect 1013 98 1014 106
rect 1016 98 1017 106
rect 1029 98 1030 106
rect 1032 98 1033 106
rect 1045 90 1046 106
rect 1048 98 1049 106
rect 1053 98 1054 106
rect 1048 90 1054 98
rect 1056 90 1057 106
rect 1061 90 1062 106
rect 1064 98 1070 106
rect 1064 90 1065 98
rect 1069 90 1070 98
rect 1072 90 1073 106
rect 1082 104 1089 106
rect 1082 100 1083 104
rect 1087 100 1089 104
rect 1082 98 1089 100
rect 1091 104 1097 106
rect 1091 100 1092 104
rect 1096 100 1097 104
rect 1091 98 1097 100
rect 1099 104 1106 106
rect 1099 100 1101 104
rect 1105 100 1106 104
rect 1099 98 1106 100
rect 1114 98 1115 106
rect 1117 98 1118 106
rect 1140 98 1142 106
rect 1144 98 1150 106
rect 1152 98 1153 106
rect 1166 98 1168 106
rect 1170 98 1172 106
rect 1467 98 1468 106
rect 1470 98 1471 106
rect 1483 98 1484 106
rect 1486 98 1487 106
rect 1499 90 1500 106
rect 1502 98 1503 106
rect 1507 98 1508 106
rect 1502 90 1508 98
rect 1510 90 1511 106
rect 1515 90 1516 106
rect 1518 98 1524 106
rect 1518 90 1519 98
rect 1523 90 1524 98
rect 1526 90 1527 106
rect 1536 104 1543 106
rect 1536 100 1537 104
rect 1541 100 1543 104
rect 1536 98 1543 100
rect 1545 104 1551 106
rect 1545 100 1546 104
rect 1550 100 1551 104
rect 1545 98 1551 100
rect 1553 104 1560 106
rect 1553 100 1555 104
rect 1559 100 1560 104
rect 1553 98 1560 100
rect 1568 98 1569 106
rect 1571 98 1572 106
rect 1596 98 1597 106
rect 1599 98 1600 106
rect 1612 98 1613 106
rect 1615 98 1616 106
rect 1628 90 1629 106
rect 1631 98 1632 106
rect 1636 98 1637 106
rect 1631 90 1637 98
rect 1639 90 1640 106
rect 1644 90 1645 106
rect 1647 98 1653 106
rect 1647 90 1648 98
rect 1652 90 1653 98
rect 1655 90 1656 106
rect 1665 104 1672 106
rect 1665 100 1666 104
rect 1670 100 1672 104
rect 1665 98 1672 100
rect 1674 104 1680 106
rect 1674 100 1675 104
rect 1679 100 1680 104
rect 1674 98 1680 100
rect 1682 104 1689 106
rect 1682 100 1684 104
rect 1688 100 1689 104
rect 1682 98 1689 100
rect 1697 98 1698 106
rect 1700 98 1701 106
rect 1723 98 1725 106
rect 1727 98 1733 106
rect 1735 98 1736 106
rect 1749 98 1751 106
rect 1753 98 1755 106
rect 9 -108 10 -100
rect 12 -108 13 -100
rect 28 -108 29 -100
rect 31 -108 32 -100
rect 50 -116 51 -100
rect 53 -116 54 -100
rect 72 -108 73 -100
rect 75 -108 76 -100
rect 88 -108 89 -100
rect 91 -108 92 -100
rect 124 -108 125 -100
rect 127 -108 128 -100
rect 146 -116 147 -100
rect 149 -116 150 -100
rect 168 -108 169 -100
rect 171 -108 172 -100
rect 184 -108 185 -100
rect 187 -108 188 -100
rect 215 -108 216 -100
rect 218 -108 219 -100
rect 255 -108 256 -100
rect 258 -108 259 -100
rect 274 -108 275 -100
rect 277 -108 278 -100
rect 296 -116 297 -100
rect 299 -116 300 -100
rect 318 -108 319 -100
rect 321 -108 322 -100
rect 334 -108 335 -100
rect 337 -108 338 -100
rect 370 -108 371 -100
rect 373 -108 374 -100
rect 392 -116 393 -100
rect 395 -116 396 -100
rect 414 -108 415 -100
rect 417 -108 418 -100
rect 430 -108 431 -100
rect 433 -108 434 -100
rect 461 -108 462 -100
rect 464 -108 465 -100
rect 756 -108 757 -100
rect 759 -108 760 -100
rect 775 -108 776 -100
rect 778 -108 779 -100
rect 797 -116 798 -100
rect 800 -116 801 -100
rect 819 -108 820 -100
rect 822 -108 823 -100
rect 835 -108 836 -100
rect 838 -108 839 -100
rect 871 -108 872 -100
rect 874 -108 875 -100
rect 893 -116 894 -100
rect 896 -116 897 -100
rect 915 -108 916 -100
rect 918 -108 919 -100
rect 931 -108 932 -100
rect 934 -108 935 -100
rect 962 -108 963 -100
rect 965 -108 966 -100
rect 1068 -108 1069 -100
rect 1071 -108 1072 -100
rect 1087 -108 1088 -100
rect 1090 -108 1091 -100
rect 1109 -116 1110 -100
rect 1112 -116 1113 -100
rect 1131 -108 1132 -100
rect 1134 -108 1135 -100
rect 1147 -108 1148 -100
rect 1150 -108 1151 -100
rect 1183 -108 1184 -100
rect 1186 -108 1187 -100
rect 1205 -116 1206 -100
rect 1208 -116 1209 -100
rect 1227 -108 1228 -100
rect 1230 -108 1231 -100
rect 1243 -108 1244 -100
rect 1246 -108 1247 -100
rect 1274 -108 1275 -100
rect 1277 -108 1278 -100
rect 1367 -108 1368 -100
rect 1370 -108 1371 -100
rect 1386 -108 1387 -100
rect 1389 -108 1390 -100
rect 1408 -116 1409 -100
rect 1411 -116 1412 -100
rect 1430 -108 1431 -100
rect 1433 -108 1434 -100
rect 1446 -108 1447 -100
rect 1449 -108 1450 -100
rect 1482 -108 1483 -100
rect 1485 -108 1486 -100
rect 1504 -116 1505 -100
rect 1507 -116 1508 -100
rect 1526 -108 1527 -100
rect 1529 -108 1530 -100
rect 1542 -108 1543 -100
rect 1545 -108 1546 -100
rect 1573 -108 1574 -100
rect 1576 -108 1577 -100
<< metal1 >>
rect -538 303 -486 307
rect -482 303 -330 307
rect -326 303 -255 307
rect -251 303 -99 307
rect -95 303 40 307
rect 44 303 196 307
rect 200 303 378 307
rect 382 303 534 307
rect 538 303 631 307
rect 635 303 787 307
rect 791 303 895 307
rect 899 303 1051 307
rect 1055 303 1179 307
rect 1183 303 1335 307
rect 1339 303 1431 307
rect 1435 303 1587 307
rect 1591 303 1690 307
rect 1694 303 1846 307
rect -538 249 -534 303
rect -514 294 -426 298
rect -422 294 -390 298
rect -386 294 -195 298
rect -191 294 -159 298
rect -155 294 100 298
rect 104 294 136 298
rect 140 294 438 298
rect 442 294 474 298
rect 478 294 691 298
rect 695 294 727 298
rect 731 294 955 298
rect 959 294 991 298
rect 995 294 1239 298
rect 1243 294 1275 298
rect 1279 294 1491 298
rect 1495 294 1527 298
rect 1531 294 1750 298
rect 1754 294 1786 298
rect -528 281 1952 282
rect -528 277 -527 281
rect -523 277 -508 281
rect -504 277 -467 281
rect -463 277 -445 281
rect -441 277 -371 281
rect -367 277 -349 281
rect -345 277 -302 281
rect -298 277 -277 281
rect -273 277 -236 281
rect -232 277 -214 281
rect -210 277 -140 281
rect -136 277 -118 281
rect -114 277 -71 281
rect -67 277 18 281
rect 22 277 59 281
rect 63 277 81 281
rect 85 277 155 281
rect 159 277 177 281
rect 181 277 224 281
rect 228 277 356 281
rect 360 277 397 281
rect 401 277 419 281
rect 423 277 493 281
rect 497 277 515 281
rect 519 277 562 281
rect 566 277 609 281
rect 613 277 650 281
rect 654 277 672 281
rect 676 277 746 281
rect 750 277 768 281
rect 772 277 815 281
rect 819 277 873 281
rect 877 277 914 281
rect 918 277 936 281
rect 940 277 1010 281
rect 1014 277 1032 281
rect 1036 277 1079 281
rect 1083 277 1157 281
rect 1161 277 1198 281
rect 1202 277 1220 281
rect 1224 277 1294 281
rect 1298 277 1316 281
rect 1320 277 1363 281
rect 1367 277 1409 281
rect 1413 277 1450 281
rect 1454 277 1472 281
rect 1476 277 1546 281
rect 1550 277 1568 281
rect 1572 277 1615 281
rect 1619 277 1668 281
rect 1672 277 1709 281
rect 1713 277 1731 281
rect 1735 277 1805 281
rect 1809 277 1827 281
rect 1831 277 1874 281
rect 1878 277 1952 281
rect -528 276 1952 277
rect -528 273 -524 276
rect -509 273 -505 276
rect -468 273 -464 276
rect -446 273 -442 276
rect -372 273 -368 276
rect -350 273 -346 276
rect -303 273 -299 276
rect -278 273 -274 276
rect -237 273 -233 276
rect -215 273 -211 276
rect -141 273 -137 276
rect -119 273 -115 276
rect -72 273 -68 276
rect 17 273 21 276
rect 58 273 62 276
rect 80 273 84 276
rect 154 273 158 276
rect 176 273 180 276
rect 223 273 227 276
rect 355 273 359 276
rect 396 273 400 276
rect 418 273 422 276
rect 492 273 496 276
rect 514 273 518 276
rect 561 273 565 276
rect 608 273 612 276
rect 649 273 653 276
rect 671 273 675 276
rect 745 273 749 276
rect 767 273 771 276
rect 814 273 818 276
rect 872 273 876 276
rect 913 273 917 276
rect 935 273 939 276
rect 1009 273 1013 276
rect 1031 273 1035 276
rect 1078 273 1082 276
rect 1156 273 1160 276
rect 1197 273 1201 276
rect 1219 273 1223 276
rect 1293 273 1297 276
rect 1315 273 1319 276
rect 1362 273 1366 276
rect 1408 273 1412 276
rect 1449 273 1453 276
rect 1471 273 1475 276
rect 1545 273 1549 276
rect 1567 273 1571 276
rect 1614 273 1618 276
rect 1667 273 1671 276
rect 1708 273 1712 276
rect 1730 273 1734 276
rect 1804 273 1808 276
rect 1826 273 1830 276
rect 1873 273 1877 276
rect -520 250 -516 265
rect -538 245 -527 249
rect -501 249 -497 265
rect -490 249 -486 265
rect -501 245 -486 249
rect -538 184 -534 245
rect -520 230 -516 245
rect -501 230 -497 245
rect -490 230 -486 245
rect -482 250 -478 265
rect -460 249 -456 257
rect -438 249 -434 265
rect -430 249 -426 265
rect -477 245 -467 249
rect -460 245 -453 249
rect -449 245 -445 249
rect -438 245 -426 249
rect -482 230 -478 245
rect -460 234 -456 245
rect -438 230 -434 245
rect -430 230 -426 245
rect -422 250 -418 265
rect -394 250 -390 265
rect -422 230 -418 245
rect -394 230 -390 245
rect -386 249 -382 265
rect -386 245 -378 249
rect -364 249 -360 257
rect -373 245 -371 249
rect -364 245 -357 249
rect -342 249 -338 265
rect -334 249 -330 265
rect -352 245 -349 249
rect -342 245 -330 249
rect -386 230 -382 245
rect -364 234 -360 245
rect -342 230 -338 245
rect -334 230 -330 245
rect -326 250 -322 265
rect -295 249 -291 265
rect -270 249 -266 265
rect -259 249 -255 265
rect -307 245 -302 249
rect -295 245 -287 249
rect -326 230 -322 245
rect -295 230 -291 245
rect -270 245 -255 249
rect -270 230 -266 245
rect -259 230 -255 245
rect -251 250 -247 265
rect -229 249 -225 257
rect -207 249 -203 265
rect -199 249 -195 265
rect -246 245 -236 249
rect -229 245 -222 249
rect -218 245 -214 249
rect -207 245 -195 249
rect -251 230 -247 245
rect -229 234 -225 245
rect -207 230 -203 245
rect -199 230 -195 245
rect -191 250 -187 265
rect -163 250 -159 265
rect -191 230 -187 245
rect -163 230 -159 245
rect -155 249 -151 265
rect -155 245 -147 249
rect -133 249 -129 257
rect -142 245 -140 249
rect -133 245 -126 249
rect -111 249 -107 265
rect -103 249 -99 265
rect -121 245 -118 249
rect -111 245 -99 249
rect -155 230 -151 245
rect -133 234 -129 245
rect -111 230 -107 245
rect -103 230 -99 245
rect -95 250 -91 265
rect -64 250 -60 265
rect -76 245 -71 249
rect -64 246 -53 250
rect -95 230 -91 245
rect -64 230 -60 246
rect 25 249 29 265
rect 36 249 40 265
rect 25 245 40 249
rect 25 230 29 245
rect 36 230 40 245
rect 44 250 48 265
rect 66 249 70 257
rect 88 249 92 265
rect 96 249 100 265
rect 49 245 59 249
rect 66 245 73 249
rect 77 245 81 249
rect 88 245 100 249
rect 44 230 48 245
rect 66 234 70 245
rect 88 230 92 245
rect 96 230 100 245
rect 104 250 108 265
rect 132 250 136 265
rect 104 230 108 245
rect 132 230 136 245
rect 140 249 144 265
rect 140 245 148 249
rect 162 249 166 257
rect 153 245 155 249
rect 162 245 169 249
rect 184 249 188 265
rect 192 249 196 265
rect 174 245 177 249
rect 184 245 196 249
rect 140 230 144 245
rect 162 234 166 245
rect 184 230 188 245
rect 192 230 196 245
rect 200 250 204 265
rect 231 250 235 265
rect 219 245 224 249
rect 231 246 239 250
rect 200 230 204 245
rect 231 230 235 246
rect 363 249 367 265
rect 374 249 378 265
rect 363 245 378 249
rect 363 230 367 245
rect 374 230 378 245
rect 382 250 386 265
rect 404 249 408 257
rect 426 249 430 265
rect 434 249 438 265
rect 387 245 397 249
rect 404 245 411 249
rect 415 245 419 249
rect 426 245 438 249
rect 382 230 386 245
rect 404 234 408 245
rect 426 230 430 245
rect 434 230 438 245
rect 442 250 446 265
rect 470 250 474 265
rect 442 230 446 245
rect 470 230 474 245
rect 478 249 482 265
rect 478 245 486 249
rect 500 249 504 257
rect 491 245 493 249
rect 500 245 507 249
rect 522 249 526 265
rect 530 249 534 265
rect 512 245 515 249
rect 522 245 534 249
rect 478 230 482 245
rect 500 234 504 245
rect 522 230 526 245
rect 530 230 534 245
rect 538 250 542 265
rect 569 250 573 265
rect 557 245 562 249
rect 569 246 577 250
rect 538 230 542 245
rect 569 230 573 246
rect 616 249 620 265
rect 627 249 631 265
rect 616 245 631 249
rect 616 230 620 245
rect 627 230 631 245
rect 635 250 639 265
rect 657 249 661 257
rect 679 249 683 265
rect 687 249 691 265
rect 640 245 650 249
rect 657 245 664 249
rect 668 245 672 249
rect 679 245 691 249
rect 635 230 639 245
rect 657 234 661 245
rect 679 230 683 245
rect 687 230 691 245
rect 695 250 699 265
rect 723 250 727 265
rect 695 230 699 245
rect 723 230 727 245
rect 731 249 735 265
rect 731 245 739 249
rect 753 249 757 257
rect 744 245 746 249
rect 753 245 760 249
rect 775 249 779 265
rect 783 249 787 265
rect 765 245 768 249
rect 775 245 787 249
rect 731 230 735 245
rect 753 234 757 245
rect 775 230 779 245
rect 783 230 787 245
rect 791 250 795 265
rect 822 250 826 265
rect 810 245 815 249
rect 822 246 834 250
rect 791 230 795 245
rect 822 230 826 246
rect 880 249 884 265
rect 891 249 895 265
rect 880 245 895 249
rect 880 230 884 245
rect 891 230 895 245
rect 899 250 903 265
rect 921 249 925 257
rect 943 249 947 265
rect 951 249 955 265
rect 904 245 914 249
rect 921 245 928 249
rect 932 245 936 249
rect 943 245 955 249
rect 899 230 903 245
rect 921 234 925 245
rect 943 230 947 245
rect 951 230 955 245
rect 959 250 963 265
rect 987 250 991 265
rect 959 230 963 245
rect 987 230 991 245
rect 995 249 999 265
rect 995 245 1003 249
rect 1017 249 1021 257
rect 1008 245 1010 249
rect 1017 245 1024 249
rect 1039 249 1043 265
rect 1047 249 1051 265
rect 1029 245 1032 249
rect 1039 245 1051 249
rect 995 230 999 245
rect 1017 234 1021 245
rect 1039 230 1043 245
rect 1047 230 1051 245
rect 1055 250 1059 265
rect 1086 250 1090 265
rect 1074 245 1079 249
rect 1086 246 1104 250
rect 1055 230 1059 245
rect 1086 230 1090 246
rect 1164 249 1168 265
rect 1175 249 1179 265
rect 1164 245 1179 249
rect 1164 230 1168 245
rect 1175 230 1179 245
rect 1183 250 1187 265
rect 1205 249 1209 257
rect 1227 249 1231 265
rect 1235 249 1239 265
rect 1188 245 1198 249
rect 1205 245 1212 249
rect 1216 245 1220 249
rect 1227 245 1239 249
rect 1183 230 1187 245
rect 1205 234 1209 245
rect 1227 230 1231 245
rect 1235 230 1239 245
rect 1243 250 1247 265
rect 1271 250 1275 265
rect 1243 230 1247 245
rect 1271 230 1275 245
rect 1279 249 1283 265
rect 1279 245 1287 249
rect 1301 249 1305 257
rect 1292 245 1294 249
rect 1301 245 1308 249
rect 1323 249 1327 265
rect 1331 249 1335 265
rect 1313 245 1316 249
rect 1323 245 1335 249
rect 1279 230 1283 245
rect 1301 234 1305 245
rect 1323 230 1327 245
rect 1331 230 1335 245
rect 1339 250 1343 265
rect 1370 250 1374 265
rect 1358 245 1363 249
rect 1370 246 1384 250
rect 1339 230 1343 245
rect 1370 230 1374 246
rect 1416 249 1420 265
rect 1427 249 1431 265
rect 1416 245 1431 249
rect 1416 230 1420 245
rect 1427 230 1431 245
rect 1435 250 1439 265
rect 1457 249 1461 257
rect 1479 249 1483 265
rect 1487 249 1491 265
rect 1440 245 1450 249
rect 1457 245 1464 249
rect 1468 245 1472 249
rect 1479 245 1491 249
rect 1435 230 1439 245
rect 1457 234 1461 245
rect 1479 230 1483 245
rect 1487 230 1491 245
rect 1495 250 1499 265
rect 1523 250 1527 265
rect 1495 230 1499 245
rect 1523 230 1527 245
rect 1531 249 1535 265
rect 1531 245 1539 249
rect 1553 249 1557 257
rect 1544 245 1546 249
rect 1553 245 1560 249
rect 1575 249 1579 265
rect 1583 249 1587 265
rect 1565 245 1568 249
rect 1575 245 1587 249
rect 1531 230 1535 245
rect 1553 234 1557 245
rect 1575 230 1579 245
rect 1583 230 1587 245
rect 1591 250 1595 265
rect 1622 250 1626 265
rect 1610 245 1615 249
rect 1622 246 1636 250
rect 1591 230 1595 245
rect 1622 230 1626 246
rect 1675 249 1679 265
rect 1686 249 1690 265
rect 1675 245 1690 249
rect 1675 230 1679 245
rect 1686 230 1690 245
rect 1694 250 1698 265
rect 1716 249 1720 257
rect 1738 249 1742 265
rect 1746 249 1750 265
rect 1699 245 1709 249
rect 1716 245 1723 249
rect 1727 245 1731 249
rect 1738 245 1750 249
rect 1694 230 1698 245
rect 1716 234 1720 245
rect 1738 230 1742 245
rect 1746 230 1750 245
rect 1754 250 1758 265
rect 1782 250 1786 265
rect 1754 230 1758 245
rect 1782 230 1786 245
rect 1790 249 1794 265
rect 1790 245 1798 249
rect 1812 249 1816 257
rect 1803 245 1805 249
rect 1812 245 1819 249
rect 1834 249 1838 265
rect 1842 249 1846 265
rect 1824 245 1827 249
rect 1834 245 1846 249
rect 1790 230 1794 245
rect 1812 234 1816 245
rect 1834 230 1838 245
rect 1842 230 1846 245
rect 1850 250 1854 265
rect 1881 250 1885 265
rect 1869 245 1874 249
rect 1881 246 1891 250
rect 1850 230 1854 245
rect 1881 230 1885 246
rect -528 223 -524 226
rect -509 223 -505 226
rect -468 223 -464 226
rect -446 223 -442 226
rect -372 223 -368 226
rect -350 223 -346 226
rect -303 223 -299 226
rect -278 223 -274 226
rect -237 223 -233 226
rect -215 223 -211 226
rect -141 223 -137 226
rect -119 223 -115 226
rect -72 223 -68 226
rect 17 223 21 226
rect 58 223 62 226
rect 80 223 84 226
rect 154 223 158 226
rect 176 223 180 226
rect 223 223 227 226
rect 355 223 359 226
rect 396 223 400 226
rect 418 223 422 226
rect 492 223 496 226
rect 514 223 518 226
rect 561 223 565 226
rect 608 223 612 226
rect 649 223 653 226
rect 671 223 675 226
rect 745 223 749 226
rect 767 223 771 226
rect 814 223 818 226
rect 872 223 876 226
rect 913 223 917 226
rect 935 223 939 226
rect 1009 223 1013 226
rect 1031 223 1035 226
rect 1078 223 1082 226
rect 1156 223 1160 226
rect 1197 223 1201 226
rect 1219 223 1223 226
rect 1293 223 1297 226
rect 1315 223 1319 226
rect 1362 223 1366 226
rect 1408 223 1412 226
rect 1449 223 1453 226
rect 1471 223 1475 226
rect 1545 223 1549 226
rect 1567 223 1571 226
rect 1614 223 1618 226
rect 1667 223 1671 226
rect 1708 223 1712 226
rect 1730 223 1734 226
rect 1804 223 1808 226
rect 1826 223 1830 226
rect 1873 223 1877 226
rect -528 222 1933 223
rect -528 218 -527 222
rect -523 218 -508 222
rect -504 218 -467 222
rect -463 218 -445 222
rect -441 218 -371 222
rect -367 218 -349 222
rect -345 218 -302 222
rect -298 218 -277 222
rect -273 218 -236 222
rect -232 218 -214 222
rect -210 218 -140 222
rect -136 218 -118 222
rect -114 218 -71 222
rect -67 218 18 222
rect 22 218 59 222
rect 63 218 81 222
rect 85 218 155 222
rect 159 218 177 222
rect 181 218 224 222
rect 228 218 356 222
rect 360 218 397 222
rect 401 218 419 222
rect 423 218 493 222
rect 497 218 515 222
rect 519 218 562 222
rect 566 218 609 222
rect 613 218 650 222
rect 654 218 672 222
rect 676 218 746 222
rect 750 218 768 222
rect 772 218 815 222
rect 819 218 873 222
rect 877 218 914 222
rect 918 218 936 222
rect 940 218 1010 222
rect 1014 218 1032 222
rect 1036 218 1079 222
rect 1083 218 1157 222
rect 1161 218 1198 222
rect 1202 218 1220 222
rect 1224 218 1294 222
rect 1298 218 1316 222
rect 1320 218 1363 222
rect 1367 218 1409 222
rect 1413 218 1450 222
rect 1454 218 1472 222
rect 1476 218 1546 222
rect 1550 218 1568 222
rect 1572 218 1615 222
rect 1619 218 1668 222
rect 1672 218 1709 222
rect 1713 218 1731 222
rect 1735 218 1805 222
rect 1809 218 1827 222
rect 1831 218 1874 222
rect 1878 218 1933 222
rect -528 217 1933 218
rect -514 189 -486 193
rect -482 189 -330 193
rect -326 189 -255 193
rect -251 189 -99 193
rect -95 189 40 193
rect 44 189 196 193
rect 200 189 378 193
rect 382 189 534 193
rect 538 189 631 193
rect 635 189 787 193
rect 791 189 895 193
rect 899 189 1051 193
rect 1055 189 1179 193
rect 1183 189 1335 193
rect 1339 189 1431 193
rect 1435 189 1587 193
rect 1591 189 1690 193
rect 1694 189 1846 193
rect -538 180 -426 184
rect -422 180 -390 184
rect -386 180 -195 184
rect -191 180 -159 184
rect -155 180 100 184
rect 104 180 136 184
rect 140 180 438 184
rect 442 180 474 184
rect 478 180 691 184
rect 695 180 727 184
rect 731 180 955 184
rect 959 180 991 184
rect 995 180 1239 184
rect 1243 180 1275 184
rect 1279 180 1491 184
rect 1495 180 1527 184
rect 1531 180 1750 184
rect 1754 180 1786 184
rect -538 -66 -534 180
rect 150 137 154 141
rect 21 130 25 133
rect 37 129 84 133
rect 37 123 41 129
rect 9 119 37 123
rect 50 119 53 123
rect 80 122 84 129
rect 166 129 213 133
rect 166 123 170 129
rect 138 119 166 123
rect 179 119 182 123
rect 209 122 213 129
rect 320 123 324 160
rect 340 149 349 153
rect 463 135 465 139
rect 352 129 399 133
rect 352 123 356 129
rect 324 119 352 123
rect 365 119 368 123
rect 395 122 399 129
rect 481 129 528 133
rect 481 123 485 129
rect 453 119 481 123
rect 494 119 497 123
rect 524 122 528 129
rect 884 123 888 151
rect 900 149 904 152
rect 1026 135 1029 139
rect 916 129 963 133
rect 916 123 920 129
rect 888 119 916 123
rect 929 119 932 123
rect 959 122 963 129
rect 1045 129 1092 133
rect 1045 123 1049 129
rect 1017 119 1045 123
rect 1058 119 1061 123
rect 1088 122 1092 129
rect 1467 123 1471 160
rect 1483 148 1487 150
rect 1610 135 1612 139
rect 1499 129 1546 133
rect 1499 123 1503 129
rect 1471 119 1499 123
rect 1512 119 1515 123
rect 1542 122 1546 129
rect 1628 129 1675 133
rect 1628 123 1632 129
rect 1600 119 1628 123
rect 1641 119 1644 123
rect 1671 122 1675 129
rect 1 114 1770 115
rect 1 110 15 114
rect 19 110 76 114
rect 80 110 93 114
rect 97 110 143 114
rect 147 110 205 114
rect 209 110 222 114
rect 226 110 258 114
rect 262 110 283 114
rect 287 110 330 114
rect 334 110 391 114
rect 395 110 408 114
rect 412 110 460 114
rect 464 110 520 114
rect 524 110 537 114
rect 541 110 573 114
rect 577 110 598 114
rect 602 110 895 114
rect 899 110 955 114
rect 959 110 972 114
rect 976 110 1024 114
rect 1028 110 1084 114
rect 1088 110 1101 114
rect 1105 110 1137 114
rect 1141 110 1162 114
rect 1166 110 1477 114
rect 1481 110 1538 114
rect 1542 110 1555 114
rect 1559 110 1607 114
rect 1611 110 1667 114
rect 1671 110 1684 114
rect 1688 110 1720 114
rect 1724 110 1745 114
rect 1749 110 1770 114
rect 1 109 1770 110
rect 1 106 5 109
rect 17 106 21 109
rect 41 106 45 109
rect -1 87 2 91
rect 9 70 13 98
rect 25 70 29 98
rect 37 90 49 94
rect 53 102 65 106
rect 75 104 79 109
rect 93 104 97 109
rect 102 106 106 109
rect 130 106 134 109
rect 146 106 150 109
rect 170 106 174 109
rect 57 76 61 90
rect 49 72 69 76
rect 9 38 13 65
rect 25 38 29 65
rect 49 42 53 72
rect 84 67 88 100
rect 110 67 114 98
rect 129 86 131 90
rect 138 70 142 98
rect 154 70 158 98
rect 166 90 178 94
rect 182 102 194 106
rect 204 104 208 109
rect 222 104 226 109
rect 231 106 235 109
rect 257 106 261 109
rect 283 106 287 109
rect 316 106 320 109
rect 332 106 336 109
rect 356 106 360 109
rect 186 76 190 90
rect 178 72 198 76
rect 84 63 103 67
rect 110 63 117 67
rect 94 42 98 63
rect 1 31 5 34
rect 17 31 21 34
rect 33 31 37 34
rect 65 31 69 34
rect 110 38 114 63
rect 138 38 142 65
rect 154 38 158 65
rect 178 42 182 72
rect 213 67 217 100
rect 239 67 243 98
rect 274 93 278 98
rect 293 93 297 98
rect 266 89 285 93
rect 293 89 301 93
rect 213 63 232 67
rect 239 63 259 67
rect 223 42 227 63
rect 74 31 78 34
rect 102 31 106 34
rect 130 31 134 34
rect 146 31 150 34
rect 162 31 166 34
rect 194 31 198 34
rect 239 38 243 63
rect 266 43 270 89
rect 293 38 297 89
rect 324 70 328 98
rect 340 70 344 98
rect 352 90 364 94
rect 368 102 380 106
rect 390 104 394 109
rect 408 104 412 109
rect 417 106 421 109
rect 445 106 449 109
rect 461 106 465 109
rect 485 106 489 109
rect 372 76 376 90
rect 364 72 384 76
rect 324 38 328 65
rect 340 38 344 65
rect 364 42 368 72
rect 399 67 403 100
rect 425 67 429 98
rect 444 86 446 90
rect 453 70 457 98
rect 469 70 473 98
rect 481 90 493 94
rect 497 102 509 106
rect 519 104 523 109
rect 537 104 541 109
rect 546 106 550 109
rect 572 106 576 109
rect 598 106 602 109
rect 880 106 884 109
rect 896 106 900 109
rect 920 106 924 109
rect 501 76 505 90
rect 493 72 513 76
rect 399 63 418 67
rect 425 63 432 67
rect 409 42 413 63
rect 203 31 207 34
rect 231 31 235 34
rect 257 31 261 35
rect 274 31 278 35
rect 283 31 287 34
rect 316 31 320 34
rect 332 31 336 34
rect 348 31 352 34
rect 380 31 384 34
rect 425 38 429 63
rect 453 38 457 65
rect 469 38 473 65
rect 493 42 497 72
rect 528 67 532 100
rect 554 67 558 98
rect 589 93 593 98
rect 608 93 612 98
rect 581 89 600 93
rect 608 89 616 93
rect 528 63 547 67
rect 554 63 574 67
rect 538 42 542 63
rect 389 31 393 34
rect 417 31 421 34
rect 445 31 449 34
rect 461 31 465 34
rect 477 31 481 34
rect 509 31 513 34
rect 554 38 558 63
rect 581 43 585 89
rect 608 38 612 89
rect 888 70 892 98
rect 904 70 908 98
rect 916 90 928 94
rect 932 102 944 106
rect 954 104 958 109
rect 972 104 976 109
rect 981 106 985 109
rect 1009 106 1013 109
rect 1025 106 1029 109
rect 1049 106 1053 109
rect 936 76 940 90
rect 928 72 948 76
rect 888 38 892 65
rect 904 38 908 65
rect 928 42 932 72
rect 963 67 967 100
rect 989 67 993 98
rect 1008 86 1010 90
rect 1017 70 1021 98
rect 1033 70 1037 98
rect 1045 90 1057 94
rect 1061 102 1073 106
rect 1083 104 1087 109
rect 1101 104 1105 109
rect 1110 106 1114 109
rect 1136 106 1140 109
rect 1162 106 1166 109
rect 1463 106 1467 109
rect 1479 106 1483 109
rect 1503 106 1507 109
rect 1065 76 1069 90
rect 1057 72 1077 76
rect 963 63 982 67
rect 989 63 996 67
rect 973 42 977 63
rect 518 31 522 34
rect 546 31 550 34
rect 572 31 576 35
rect 589 31 593 35
rect 598 31 602 34
rect 880 31 884 34
rect 896 31 900 34
rect 912 31 916 34
rect 944 31 948 34
rect 989 38 993 63
rect 1017 38 1021 65
rect 1033 38 1037 65
rect 1057 42 1061 72
rect 1092 67 1096 100
rect 1118 67 1122 98
rect 1153 93 1157 98
rect 1172 93 1176 98
rect 1145 89 1164 93
rect 1172 89 1180 93
rect 1092 63 1111 67
rect 1118 63 1138 67
rect 1102 42 1106 63
rect 953 31 957 34
rect 981 31 985 34
rect 1009 31 1013 34
rect 1025 31 1029 34
rect 1041 31 1045 34
rect 1073 31 1077 34
rect 1118 38 1122 63
rect 1145 43 1149 89
rect 1172 38 1176 89
rect 1471 70 1475 98
rect 1487 70 1491 98
rect 1499 90 1511 94
rect 1515 102 1527 106
rect 1537 104 1541 109
rect 1555 104 1559 109
rect 1564 106 1568 109
rect 1592 106 1596 109
rect 1608 106 1612 109
rect 1632 106 1636 109
rect 1519 76 1523 90
rect 1511 72 1531 76
rect 1471 38 1475 65
rect 1487 38 1491 65
rect 1511 42 1515 72
rect 1546 67 1550 100
rect 1572 67 1576 98
rect 1591 86 1593 90
rect 1600 70 1604 98
rect 1616 70 1620 98
rect 1628 90 1640 94
rect 1644 102 1656 106
rect 1666 104 1670 109
rect 1684 104 1688 109
rect 1693 106 1697 109
rect 1719 106 1723 109
rect 1745 106 1749 109
rect 1648 76 1652 90
rect 1640 72 1660 76
rect 1546 63 1565 67
rect 1572 63 1579 67
rect 1556 42 1560 63
rect 1082 31 1086 34
rect 1110 31 1114 34
rect 1136 31 1140 35
rect 1153 31 1157 35
rect 1162 31 1166 34
rect 1463 31 1467 34
rect 1479 31 1483 34
rect 1495 31 1499 34
rect 1527 31 1531 34
rect 1572 38 1576 63
rect 1600 38 1604 65
rect 1616 38 1620 65
rect 1640 42 1644 72
rect 1675 67 1679 100
rect 1701 67 1705 98
rect 1736 93 1740 98
rect 1755 93 1759 98
rect 1728 89 1747 93
rect 1755 89 1806 93
rect 1675 63 1694 67
rect 1701 63 1721 67
rect 1685 42 1689 63
rect 1536 31 1540 34
rect 1564 31 1568 34
rect 1592 31 1596 34
rect 1608 31 1612 34
rect 1624 31 1628 34
rect 1656 31 1660 34
rect 1701 38 1705 63
rect 1728 43 1732 89
rect 1755 38 1759 89
rect 1802 59 1806 89
rect 1665 31 1669 34
rect 1693 31 1697 34
rect 1719 31 1723 35
rect 1736 31 1740 35
rect 1745 31 1749 34
rect 1927 31 1933 217
rect 0 30 1933 31
rect 0 26 2 30
rect 6 26 75 30
rect 79 26 93 30
rect 97 26 103 30
rect 107 26 131 30
rect 135 26 204 30
rect 208 26 222 30
rect 226 26 232 30
rect 236 26 265 30
rect 269 26 283 30
rect 287 26 317 30
rect 321 26 390 30
rect 394 26 408 30
rect 412 26 418 30
rect 422 26 446 30
rect 450 26 519 30
rect 523 26 537 30
rect 541 26 547 30
rect 551 26 580 30
rect 584 26 598 30
rect 602 26 881 30
rect 885 26 954 30
rect 958 26 972 30
rect 976 26 982 30
rect 986 26 1010 30
rect 1014 26 1083 30
rect 1087 26 1101 30
rect 1105 26 1111 30
rect 1115 26 1144 30
rect 1148 26 1162 30
rect 1166 26 1464 30
rect 1468 26 1537 30
rect 1541 26 1555 30
rect 1559 26 1565 30
rect 1569 26 1593 30
rect 1597 26 1666 30
rect 1670 26 1684 30
rect 1688 26 1694 30
rect 1698 26 1727 30
rect 1731 26 1745 30
rect 1749 26 1933 30
rect 0 25 1933 26
rect 25 17 45 21
rect 45 10 49 17
rect 58 17 61 21
rect 88 10 92 18
rect 154 17 174 21
rect 45 6 92 10
rect 174 10 178 17
rect 187 17 190 21
rect 217 10 221 18
rect 270 16 274 18
rect 340 17 360 21
rect 174 6 221 10
rect 360 10 364 17
rect 373 17 376 21
rect 403 10 407 18
rect 469 17 489 21
rect 360 6 407 10
rect 489 10 493 17
rect 502 17 505 21
rect 532 10 536 18
rect 585 16 589 18
rect 904 17 924 21
rect 489 6 536 10
rect 924 10 928 17
rect 937 17 940 21
rect 967 10 971 18
rect 1033 17 1053 21
rect 924 6 971 10
rect 1053 10 1057 17
rect 1066 17 1069 21
rect 1096 10 1100 18
rect 1149 16 1153 18
rect 1487 17 1507 21
rect 1053 6 1100 10
rect 1507 10 1511 17
rect 1520 17 1523 21
rect 1550 10 1554 18
rect 1616 17 1636 21
rect 1507 6 1554 10
rect 1636 10 1640 17
rect 1649 17 1652 21
rect 1679 10 1683 18
rect 1732 16 1736 18
rect 1636 6 1683 10
rect 1802 -35 1806 -3
rect 1344 -39 1806 -35
rect 9 -53 13 -49
rect -538 -70 28 -66
rect 32 -70 184 -66
rect 188 -70 274 -66
rect 278 -70 430 -66
rect 434 -70 775 -66
rect 779 -70 931 -66
rect 935 -70 1087 -66
rect 1091 -70 1243 -66
rect 1247 -70 1386 -66
rect 1390 -70 1542 -66
rect -538 -189 -534 -70
rect -4 -79 88 -75
rect 92 -79 124 -75
rect 128 -79 334 -75
rect 338 -79 370 -75
rect 374 -79 835 -75
rect 839 -79 871 -75
rect 875 -79 1147 -75
rect 1151 -79 1183 -75
rect 1187 -79 1446 -75
rect 1450 -79 1482 -75
rect 3 -92 1581 -91
rect 3 -96 4 -92
rect 8 -96 47 -92
rect 51 -96 69 -92
rect 73 -96 143 -92
rect 147 -96 165 -92
rect 169 -96 212 -92
rect 216 -96 252 -92
rect 256 -96 293 -92
rect 297 -96 315 -92
rect 319 -96 389 -92
rect 393 -96 411 -92
rect 415 -96 458 -92
rect 462 -96 753 -92
rect 757 -96 794 -92
rect 798 -96 816 -92
rect 820 -96 890 -92
rect 894 -96 912 -92
rect 916 -96 959 -92
rect 963 -96 1065 -92
rect 1069 -96 1106 -92
rect 1110 -96 1128 -92
rect 1132 -96 1202 -92
rect 1206 -96 1224 -92
rect 1228 -96 1271 -92
rect 1275 -96 1364 -92
rect 1368 -96 1405 -92
rect 1409 -96 1427 -92
rect 1431 -96 1501 -92
rect 1505 -96 1523 -92
rect 1527 -96 1570 -92
rect 1574 -96 1581 -92
rect 3 -97 1581 -96
rect 5 -100 9 -97
rect 46 -100 50 -97
rect 68 -100 72 -97
rect 142 -100 146 -97
rect 164 -100 168 -97
rect 211 -100 215 -97
rect 251 -100 255 -97
rect 292 -100 296 -97
rect 314 -100 318 -97
rect 388 -100 392 -97
rect 410 -100 414 -97
rect 457 -100 461 -97
rect 752 -100 756 -97
rect 793 -100 797 -97
rect 815 -100 819 -97
rect 889 -100 893 -97
rect 911 -100 915 -97
rect 958 -100 962 -97
rect 1064 -100 1068 -97
rect 1105 -100 1109 -97
rect 1127 -100 1131 -97
rect 1201 -100 1205 -97
rect 1223 -100 1227 -97
rect 1270 -100 1274 -97
rect 1363 -100 1367 -97
rect 1404 -100 1408 -97
rect 1426 -100 1430 -97
rect 1500 -100 1504 -97
rect 1522 -100 1526 -97
rect 1569 -100 1573 -97
rect 13 -124 17 -108
rect 24 -124 28 -108
rect 13 -128 28 -124
rect 13 -143 17 -128
rect 24 -143 28 -128
rect 32 -123 36 -108
rect 54 -124 58 -116
rect 76 -124 80 -108
rect 84 -124 88 -108
rect 37 -128 47 -124
rect 54 -128 61 -124
rect 65 -128 69 -124
rect 76 -128 88 -124
rect 32 -143 36 -128
rect 54 -139 58 -128
rect 76 -143 80 -128
rect 84 -143 88 -128
rect 92 -123 96 -108
rect 120 -123 124 -108
rect 92 -143 96 -128
rect 120 -143 124 -128
rect 128 -124 132 -108
rect 128 -128 136 -124
rect 150 -124 154 -116
rect 141 -128 143 -124
rect 150 -128 157 -124
rect 172 -124 176 -108
rect 180 -124 184 -108
rect 162 -128 165 -124
rect 172 -128 184 -124
rect 128 -143 132 -128
rect 150 -139 154 -128
rect 172 -143 176 -128
rect 180 -143 184 -128
rect 188 -123 192 -108
rect 219 -124 223 -108
rect 207 -128 212 -124
rect 219 -128 227 -124
rect 259 -124 263 -108
rect 270 -124 274 -108
rect 250 -128 252 -124
rect 259 -128 274 -124
rect 188 -143 192 -128
rect 219 -143 223 -128
rect 259 -143 263 -128
rect 270 -143 274 -128
rect 278 -123 282 -108
rect 300 -124 304 -116
rect 322 -124 326 -108
rect 330 -124 334 -108
rect 283 -128 293 -124
rect 300 -128 307 -124
rect 311 -128 315 -124
rect 322 -128 334 -124
rect 278 -143 282 -128
rect 300 -139 304 -128
rect 322 -143 326 -128
rect 330 -143 334 -128
rect 338 -123 342 -108
rect 366 -123 370 -108
rect 338 -143 342 -128
rect 366 -143 370 -128
rect 374 -124 378 -108
rect 374 -128 382 -124
rect 396 -124 400 -116
rect 387 -128 389 -124
rect 396 -128 403 -124
rect 418 -124 422 -108
rect 426 -124 430 -108
rect 408 -128 411 -124
rect 418 -128 430 -124
rect 374 -143 378 -128
rect 396 -139 400 -128
rect 418 -143 422 -128
rect 426 -143 430 -128
rect 434 -123 438 -108
rect 465 -124 469 -108
rect 453 -128 458 -124
rect 465 -128 473 -124
rect 760 -124 764 -108
rect 771 -124 775 -108
rect 744 -128 753 -124
rect 760 -128 775 -124
rect 434 -143 438 -128
rect 465 -143 469 -128
rect 760 -143 764 -128
rect 771 -143 775 -128
rect 779 -123 783 -108
rect 801 -124 805 -116
rect 823 -124 827 -108
rect 831 -124 835 -108
rect 784 -128 794 -124
rect 801 -128 808 -124
rect 812 -128 816 -124
rect 823 -128 835 -124
rect 779 -143 783 -128
rect 801 -139 805 -128
rect 823 -143 827 -128
rect 831 -143 835 -128
rect 839 -123 843 -108
rect 867 -123 871 -108
rect 839 -143 843 -128
rect 867 -143 871 -128
rect 875 -124 879 -108
rect 875 -128 883 -124
rect 897 -124 901 -116
rect 888 -128 890 -124
rect 897 -128 904 -124
rect 919 -124 923 -108
rect 927 -124 931 -108
rect 909 -128 912 -124
rect 919 -128 931 -124
rect 875 -143 879 -128
rect 897 -139 901 -128
rect 919 -143 923 -128
rect 927 -143 931 -128
rect 935 -123 939 -108
rect 966 -124 970 -108
rect 954 -128 959 -124
rect 966 -128 974 -124
rect 1072 -124 1076 -108
rect 1083 -124 1087 -108
rect 1047 -128 1065 -124
rect 1072 -128 1087 -124
rect 935 -143 939 -128
rect 966 -143 970 -128
rect 1072 -143 1076 -128
rect 1083 -143 1087 -128
rect 1091 -123 1095 -108
rect 1113 -124 1117 -116
rect 1135 -124 1139 -108
rect 1143 -124 1147 -108
rect 1096 -128 1106 -124
rect 1113 -128 1120 -124
rect 1124 -128 1128 -124
rect 1135 -128 1147 -124
rect 1091 -143 1095 -128
rect 1113 -139 1117 -128
rect 1135 -143 1139 -128
rect 1143 -143 1147 -128
rect 1151 -123 1155 -108
rect 1179 -123 1183 -108
rect 1151 -143 1155 -128
rect 1179 -143 1183 -128
rect 1187 -124 1191 -108
rect 1187 -128 1195 -124
rect 1209 -124 1213 -116
rect 1200 -128 1202 -124
rect 1209 -128 1216 -124
rect 1231 -124 1235 -108
rect 1239 -124 1243 -108
rect 1221 -128 1224 -124
rect 1231 -128 1243 -124
rect 1187 -143 1191 -128
rect 1209 -139 1213 -128
rect 1231 -143 1235 -128
rect 1239 -143 1243 -128
rect 1247 -123 1251 -108
rect 1278 -124 1282 -108
rect 1266 -128 1271 -124
rect 1278 -128 1286 -124
rect 1371 -124 1375 -108
rect 1382 -124 1386 -108
rect 1344 -128 1364 -124
rect 1371 -128 1386 -124
rect 1247 -143 1251 -128
rect 1278 -143 1282 -128
rect 1371 -143 1375 -128
rect 1382 -143 1386 -128
rect 1390 -123 1394 -108
rect 1412 -124 1416 -116
rect 1434 -124 1438 -108
rect 1442 -124 1446 -108
rect 1395 -128 1405 -124
rect 1412 -128 1419 -124
rect 1423 -128 1427 -124
rect 1434 -128 1446 -124
rect 1390 -143 1394 -128
rect 1412 -139 1416 -128
rect 1434 -143 1438 -128
rect 1442 -143 1446 -128
rect 1450 -123 1454 -108
rect 1478 -123 1482 -108
rect 1450 -143 1454 -128
rect 1478 -143 1482 -128
rect 1486 -124 1490 -108
rect 1486 -128 1494 -124
rect 1508 -124 1512 -116
rect 1499 -128 1501 -124
rect 1508 -128 1515 -124
rect 1530 -124 1534 -108
rect 1538 -124 1542 -108
rect 1520 -128 1523 -124
rect 1530 -128 1542 -124
rect 1486 -143 1490 -128
rect 1508 -139 1512 -128
rect 1530 -143 1534 -128
rect 1538 -143 1542 -128
rect 1546 -123 1550 -108
rect 1577 -124 1581 -108
rect 1565 -128 1570 -124
rect 1577 -128 1585 -124
rect 1546 -143 1550 -128
rect 1577 -143 1581 -128
rect 5 -150 9 -147
rect 46 -150 50 -147
rect 68 -150 72 -147
rect 142 -150 146 -147
rect 164 -150 168 -147
rect 211 -150 215 -147
rect 251 -150 255 -147
rect 292 -150 296 -147
rect 314 -150 318 -147
rect 388 -150 392 -147
rect 410 -150 414 -147
rect 457 -150 461 -147
rect 752 -150 756 -147
rect 793 -150 797 -147
rect 815 -150 819 -147
rect 889 -150 893 -147
rect 911 -150 915 -147
rect 958 -150 962 -147
rect 1064 -150 1068 -147
rect 1105 -150 1109 -147
rect 1127 -150 1131 -147
rect 1201 -150 1205 -147
rect 1223 -150 1227 -147
rect 1270 -150 1274 -147
rect 1363 -150 1367 -147
rect 1404 -150 1408 -147
rect 1426 -150 1430 -147
rect 1500 -150 1504 -147
rect 1522 -150 1526 -147
rect 1569 -150 1573 -147
rect 1927 -150 1933 25
rect 3 -151 1933 -150
rect 3 -155 6 -151
rect 10 -155 47 -151
rect 51 -155 69 -151
rect 73 -155 143 -151
rect 147 -155 165 -151
rect 169 -155 212 -151
rect 216 -155 252 -151
rect 256 -155 293 -151
rect 297 -155 315 -151
rect 319 -155 389 -151
rect 393 -155 411 -151
rect 415 -155 458 -151
rect 462 -155 753 -151
rect 757 -155 794 -151
rect 798 -155 816 -151
rect 820 -155 890 -151
rect 894 -155 912 -151
rect 916 -155 959 -151
rect 963 -155 1065 -151
rect 1069 -155 1106 -151
rect 1110 -155 1128 -151
rect 1132 -155 1202 -151
rect 1206 -155 1224 -151
rect 1228 -155 1271 -151
rect 1275 -155 1364 -151
rect 1368 -155 1405 -151
rect 1409 -155 1427 -151
rect 1431 -155 1501 -151
rect 1505 -155 1523 -151
rect 1527 -155 1570 -151
rect 1574 -155 1933 -151
rect 3 -156 1933 -155
rect 3 -184 28 -180
rect 32 -184 184 -180
rect 188 -184 274 -180
rect 278 -184 430 -180
rect 434 -184 775 -180
rect 779 -184 931 -180
rect 935 -184 1087 -180
rect 1091 -184 1243 -180
rect 1247 -184 1386 -180
rect 1390 -184 1542 -180
rect 1927 -187 1933 -156
rect -538 -193 88 -189
rect 92 -193 124 -189
rect 128 -193 334 -189
rect 338 -193 370 -189
rect 374 -193 835 -189
rect 839 -193 871 -189
rect 875 -193 1147 -189
rect 1151 -193 1183 -189
rect 1187 -193 1446 -189
rect 1450 -193 1482 -189
rect -538 -205 -534 -193
<< metal2 >>
rect -486 303 -482 307
rect -255 303 -251 307
rect 40 303 44 307
rect 378 303 382 307
rect 631 303 635 307
rect 895 303 899 307
rect 1179 303 1183 307
rect 1431 303 1435 307
rect 1690 303 1694 307
rect -390 294 -386 298
rect -159 294 -155 298
rect 136 294 140 298
rect 474 294 478 298
rect 727 294 731 298
rect 991 294 995 298
rect 1275 294 1279 298
rect 1527 294 1531 298
rect 1786 294 1790 298
rect -519 250 -515 293
rect -453 285 -391 289
rect -519 194 -515 245
rect -453 249 -449 285
rect -395 250 -391 285
rect -357 285 -308 289
rect -357 250 -353 285
rect -312 250 -308 285
rect -222 285 -160 289
rect -482 223 -478 245
rect -421 223 -417 245
rect -482 219 -417 223
rect -377 216 -373 245
rect -325 216 -321 245
rect -377 212 -321 216
rect -486 189 -482 193
rect -330 189 -326 193
rect -519 -75 -515 189
rect -390 180 -386 184
rect -286 91 -282 244
rect -222 249 -218 285
rect -164 250 -160 285
rect -126 285 -77 289
rect -126 250 -122 285
rect -81 250 -77 285
rect 73 285 135 289
rect -251 223 -247 245
rect -190 223 -186 245
rect -251 219 -186 223
rect -146 216 -142 245
rect -94 216 -90 245
rect -146 212 -90 216
rect -255 189 -251 193
rect -99 189 -95 193
rect -159 180 -155 184
rect -52 148 -48 245
rect 73 249 77 285
rect 131 250 135 285
rect 169 285 218 289
rect 169 250 173 285
rect 214 250 218 285
rect 411 285 473 289
rect 44 223 48 245
rect 105 223 109 245
rect 44 219 109 223
rect 149 216 153 245
rect 201 216 205 245
rect 149 212 205 216
rect 40 189 44 193
rect 196 189 200 193
rect 136 180 140 184
rect 240 164 244 245
rect 411 249 415 285
rect 469 250 473 285
rect 507 285 556 289
rect 507 250 511 285
rect 552 250 556 285
rect 664 285 726 289
rect 382 223 386 245
rect 443 223 447 245
rect 382 219 447 223
rect 487 216 491 245
rect 539 216 543 245
rect 487 212 543 216
rect 378 189 382 193
rect 534 189 538 193
rect 474 180 478 184
rect 578 165 582 245
rect 664 249 668 285
rect 722 250 726 285
rect 760 285 809 289
rect 760 250 764 285
rect 805 250 809 285
rect 928 285 990 289
rect 635 223 639 245
rect 696 223 700 245
rect 635 219 700 223
rect 740 216 744 245
rect 792 216 796 245
rect 740 212 796 216
rect 631 189 635 193
rect 787 189 791 193
rect 727 180 731 184
rect 150 160 244 164
rect 325 161 582 165
rect -52 144 25 148
rect 150 146 154 160
rect 835 153 839 245
rect 928 249 932 285
rect 986 250 990 285
rect 1024 285 1073 289
rect 1024 250 1028 285
rect 1069 250 1073 285
rect 1212 285 1274 289
rect 899 223 903 245
rect 960 223 964 245
rect 899 219 964 223
rect 1004 216 1008 245
rect 1056 216 1060 245
rect 1004 212 1060 216
rect 895 189 899 193
rect 1051 189 1055 193
rect 991 180 995 184
rect 1105 175 1109 245
rect 1212 249 1216 285
rect 1270 250 1274 285
rect 1308 285 1357 289
rect 1308 250 1312 285
rect 1353 250 1357 285
rect 1464 285 1526 289
rect 1183 223 1187 245
rect 1244 223 1248 245
rect 1183 219 1248 223
rect 1288 216 1292 245
rect 1340 216 1344 245
rect 1288 212 1344 216
rect 1179 189 1183 193
rect 1335 189 1339 193
rect 1275 180 1279 184
rect 884 171 1109 175
rect 884 156 888 171
rect 1384 157 1389 245
rect 1464 249 1468 285
rect 1522 250 1526 285
rect 1560 285 1609 289
rect 1560 250 1564 285
rect 1605 250 1609 285
rect 1723 285 1785 289
rect 1435 223 1439 245
rect 1496 223 1500 245
rect 1435 219 1500 223
rect 1540 216 1544 245
rect 1592 216 1596 245
rect 1540 212 1596 216
rect 1431 189 1435 193
rect 1587 189 1591 193
rect 1527 180 1531 184
rect 1637 174 1641 245
rect 1723 249 1727 285
rect 1781 250 1785 285
rect 1819 285 1868 289
rect 1819 250 1823 285
rect 1864 250 1868 285
rect 1694 223 1698 245
rect 1755 223 1759 245
rect 1694 219 1759 223
rect 1799 216 1803 245
rect 1851 216 1855 245
rect 1799 212 1855 216
rect 1690 189 1694 193
rect 1846 189 1850 193
rect 1786 180 1790 184
rect 1467 170 1641 174
rect 1467 165 1472 170
rect 1892 159 1896 245
rect 354 149 839 153
rect 905 153 1389 157
rect 1482 155 1896 159
rect 21 138 25 144
rect 302 135 458 139
rect 617 135 1021 139
rect 46 115 50 119
rect 175 115 179 119
rect 26 111 50 115
rect 155 111 179 115
rect -286 87 -6 91
rect 26 70 30 111
rect 124 75 128 85
rect 74 71 128 75
rect 155 70 159 111
rect 302 94 306 135
rect 361 115 365 119
rect 490 115 494 119
rect 341 111 365 115
rect 470 111 494 115
rect 203 71 306 75
rect 10 29 14 65
rect 10 25 57 29
rect 53 21 57 25
rect 118 4 122 62
rect 139 29 143 65
rect 139 25 186 29
rect 182 21 186 25
rect 269 4 273 11
rect 118 0 273 4
rect 302 -9 306 71
rect 341 70 345 111
rect 439 75 443 85
rect 389 71 443 75
rect 470 70 474 111
rect 617 94 621 135
rect 1181 135 1605 139
rect 925 115 929 119
rect 1054 115 1058 119
rect 905 111 929 115
rect 1034 111 1058 115
rect 518 71 626 75
rect 325 29 329 65
rect 325 25 372 29
rect 368 21 372 25
rect 433 4 437 62
rect 454 29 458 65
rect 454 25 501 29
rect 497 21 501 25
rect 584 4 588 11
rect 433 0 588 4
rect 9 -13 306 -9
rect 9 -44 13 -13
rect 622 -29 626 71
rect 905 70 909 111
rect 1003 75 1007 85
rect 953 71 1007 75
rect 1034 70 1038 111
rect 1181 94 1185 135
rect 1508 115 1512 119
rect 1637 115 1641 119
rect 1488 111 1512 115
rect 1617 111 1641 115
rect 1082 71 1198 75
rect 889 29 893 65
rect 889 25 936 29
rect 932 21 936 25
rect 997 4 1001 62
rect 1018 29 1022 65
rect 1018 25 1065 29
rect 1061 21 1065 25
rect 1148 4 1152 11
rect 997 0 1152 4
rect 1194 -4 1198 71
rect 1488 70 1492 111
rect 1586 75 1590 85
rect 1536 71 1590 75
rect 1617 70 1621 111
rect 1954 115 1960 274
rect 1778 109 1960 115
rect 1665 71 1783 75
rect 1472 29 1476 65
rect 1472 25 1519 29
rect 1515 21 1519 25
rect 1580 4 1584 62
rect 1601 29 1605 65
rect 1601 25 1648 29
rect 1644 21 1648 25
rect 1731 4 1735 11
rect 1580 0 1735 4
rect 237 -33 626 -29
rect 739 -8 1198 -4
rect 28 -70 32 -66
rect -519 -79 -9 -75
rect -519 -180 -515 -79
rect 124 -79 128 -75
rect 61 -88 123 -84
rect 61 -124 65 -88
rect 119 -123 123 -88
rect 157 -88 206 -84
rect 157 -123 161 -88
rect 202 -123 206 -88
rect 237 -124 241 -33
rect 274 -70 278 -66
rect 370 -79 374 -75
rect 307 -88 369 -84
rect 237 -128 245 -124
rect 307 -124 311 -88
rect 365 -123 369 -88
rect 403 -88 452 -84
rect 403 -123 407 -88
rect 448 -123 452 -88
rect 739 -123 743 -8
rect 1779 -18 1783 71
rect 1802 2 1806 54
rect 1042 -22 1783 -18
rect 775 -70 779 -66
rect 871 -79 875 -75
rect 808 -88 870 -84
rect 808 -124 812 -88
rect 866 -123 870 -88
rect 904 -88 953 -84
rect 904 -123 908 -88
rect 949 -123 953 -88
rect 1042 -123 1046 -22
rect 1087 -70 1091 -66
rect 1183 -79 1187 -75
rect 1120 -88 1182 -84
rect 1120 -124 1124 -88
rect 1178 -123 1182 -88
rect 1216 -88 1265 -84
rect 1216 -123 1220 -88
rect 1261 -123 1265 -88
rect 1339 -123 1343 -40
rect 1386 -70 1390 -66
rect 1482 -79 1486 -75
rect 1419 -88 1481 -84
rect 1419 -124 1423 -88
rect 1477 -123 1481 -88
rect 1515 -88 1564 -84
rect 1515 -123 1519 -88
rect 1560 -123 1564 -88
rect 1954 -91 1960 109
rect 1589 -97 1960 -91
rect 32 -150 36 -128
rect 93 -150 97 -128
rect 32 -154 97 -150
rect 137 -157 141 -128
rect 189 -157 193 -128
rect 278 -150 282 -128
rect 339 -150 343 -128
rect 278 -154 343 -150
rect 137 -161 193 -157
rect 383 -157 387 -128
rect 435 -157 439 -128
rect 779 -150 783 -128
rect 840 -150 844 -128
rect 779 -154 844 -150
rect 383 -161 439 -157
rect 884 -157 888 -128
rect 936 -157 940 -128
rect 1091 -150 1095 -128
rect 1152 -150 1156 -128
rect 1091 -154 1156 -150
rect 884 -161 940 -157
rect 1196 -157 1200 -128
rect 1248 -157 1252 -128
rect 1390 -150 1394 -128
rect 1451 -150 1455 -128
rect 1390 -154 1455 -150
rect 1196 -161 1252 -157
rect 1495 -157 1499 -128
rect 1547 -157 1551 -128
rect 1495 -161 1551 -157
rect -519 -184 -2 -180
rect 28 -184 32 -180
rect 184 -184 188 -180
rect 274 -184 278 -180
rect 430 -184 434 -180
rect 775 -184 779 -180
rect 931 -184 935 -180
rect 1087 -184 1091 -180
rect 1243 -184 1247 -180
rect 1386 -184 1390 -180
rect 1542 -184 1546 -180
rect -519 -204 -515 -184
rect 1954 -186 1960 -97
rect 124 -193 128 -189
rect 370 -193 374 -189
rect 871 -193 875 -189
rect 1183 -193 1187 -189
rect 1482 -193 1486 -189
<< ntransistor >>
rect -523 226 -521 230
rect -504 226 -502 230
rect -485 226 -483 230
rect -463 226 -461 234
rect -441 226 -439 230
rect -425 226 -423 230
rect -389 226 -387 230
rect -367 226 -365 234
rect -345 226 -343 230
rect -329 226 -327 230
rect -298 226 -296 230
rect -273 226 -271 230
rect -254 226 -252 230
rect -232 226 -230 234
rect -210 226 -208 230
rect -194 226 -192 230
rect -158 226 -156 230
rect -136 226 -134 234
rect -114 226 -112 230
rect -98 226 -96 230
rect -67 226 -65 230
rect 22 226 24 230
rect 41 226 43 230
rect 63 226 65 234
rect 85 226 87 230
rect 101 226 103 230
rect 137 226 139 230
rect 159 226 161 234
rect 181 226 183 230
rect 197 226 199 230
rect 228 226 230 230
rect 360 226 362 230
rect 379 226 381 230
rect 401 226 403 234
rect 423 226 425 230
rect 439 226 441 230
rect 475 226 477 230
rect 497 226 499 234
rect 519 226 521 230
rect 535 226 537 230
rect 566 226 568 230
rect 613 226 615 230
rect 632 226 634 230
rect 654 226 656 234
rect 676 226 678 230
rect 692 226 694 230
rect 728 226 730 230
rect 750 226 752 234
rect 772 226 774 230
rect 788 226 790 230
rect 819 226 821 230
rect 877 226 879 230
rect 896 226 898 230
rect 918 226 920 234
rect 940 226 942 230
rect 956 226 958 230
rect 992 226 994 230
rect 1014 226 1016 234
rect 1036 226 1038 230
rect 1052 226 1054 230
rect 1083 226 1085 230
rect 1161 226 1163 230
rect 1180 226 1182 230
rect 1202 226 1204 234
rect 1224 226 1226 230
rect 1240 226 1242 230
rect 1276 226 1278 230
rect 1298 226 1300 234
rect 1320 226 1322 230
rect 1336 226 1338 230
rect 1367 226 1369 230
rect 1413 226 1415 230
rect 1432 226 1434 230
rect 1454 226 1456 234
rect 1476 226 1478 230
rect 1492 226 1494 230
rect 1528 226 1530 230
rect 1550 226 1552 234
rect 1572 226 1574 230
rect 1588 226 1590 230
rect 1619 226 1621 230
rect 1672 226 1674 230
rect 1691 226 1693 230
rect 1713 226 1715 234
rect 1735 226 1737 230
rect 1751 226 1753 230
rect 1787 226 1789 230
rect 1809 226 1811 234
rect 1831 226 1833 230
rect 1847 226 1849 230
rect 1878 226 1880 230
rect 6 34 8 38
rect 22 34 24 38
rect 38 34 40 42
rect 46 34 48 42
rect 54 34 56 42
rect 62 34 64 42
rect 81 34 83 42
rect 89 34 91 42
rect 107 34 109 38
rect 135 34 137 38
rect 151 34 153 38
rect 167 34 169 42
rect 175 34 177 42
rect 183 34 185 42
rect 191 34 193 42
rect 210 34 212 42
rect 218 34 220 42
rect 236 34 238 38
rect 263 35 265 43
rect 271 35 273 43
rect 289 34 291 38
rect 321 34 323 38
rect 337 34 339 38
rect 353 34 355 42
rect 361 34 363 42
rect 369 34 371 42
rect 377 34 379 42
rect 396 34 398 42
rect 404 34 406 42
rect 422 34 424 38
rect 450 34 452 38
rect 466 34 468 38
rect 482 34 484 42
rect 490 34 492 42
rect 498 34 500 42
rect 506 34 508 42
rect 525 34 527 42
rect 533 34 535 42
rect 551 34 553 38
rect 578 35 580 43
rect 586 35 588 43
rect 604 34 606 38
rect 885 34 887 38
rect 901 34 903 38
rect 917 34 919 42
rect 925 34 927 42
rect 933 34 935 42
rect 941 34 943 42
rect 960 34 962 42
rect 968 34 970 42
rect 986 34 988 38
rect 1014 34 1016 38
rect 1030 34 1032 38
rect 1046 34 1048 42
rect 1054 34 1056 42
rect 1062 34 1064 42
rect 1070 34 1072 42
rect 1089 34 1091 42
rect 1097 34 1099 42
rect 1115 34 1117 38
rect 1142 35 1144 43
rect 1150 35 1152 43
rect 1168 34 1170 38
rect 1468 34 1470 38
rect 1484 34 1486 38
rect 1500 34 1502 42
rect 1508 34 1510 42
rect 1516 34 1518 42
rect 1524 34 1526 42
rect 1543 34 1545 42
rect 1551 34 1553 42
rect 1569 34 1571 38
rect 1597 34 1599 38
rect 1613 34 1615 38
rect 1629 34 1631 42
rect 1637 34 1639 42
rect 1645 34 1647 42
rect 1653 34 1655 42
rect 1672 34 1674 42
rect 1680 34 1682 42
rect 1698 34 1700 38
rect 1725 35 1727 43
rect 1733 35 1735 43
rect 1751 34 1753 38
rect 10 -147 12 -143
rect 29 -147 31 -143
rect 51 -147 53 -139
rect 73 -147 75 -143
rect 89 -147 91 -143
rect 125 -147 127 -143
rect 147 -147 149 -139
rect 169 -147 171 -143
rect 185 -147 187 -143
rect 216 -147 218 -143
rect 256 -147 258 -143
rect 275 -147 277 -143
rect 297 -147 299 -139
rect 319 -147 321 -143
rect 335 -147 337 -143
rect 371 -147 373 -143
rect 393 -147 395 -139
rect 415 -147 417 -143
rect 431 -147 433 -143
rect 462 -147 464 -143
rect 757 -147 759 -143
rect 776 -147 778 -143
rect 798 -147 800 -139
rect 820 -147 822 -143
rect 836 -147 838 -143
rect 872 -147 874 -143
rect 894 -147 896 -139
rect 916 -147 918 -143
rect 932 -147 934 -143
rect 963 -147 965 -143
rect 1069 -147 1071 -143
rect 1088 -147 1090 -143
rect 1110 -147 1112 -139
rect 1132 -147 1134 -143
rect 1148 -147 1150 -143
rect 1184 -147 1186 -143
rect 1206 -147 1208 -139
rect 1228 -147 1230 -143
rect 1244 -147 1246 -143
rect 1275 -147 1277 -143
rect 1368 -147 1370 -143
rect 1387 -147 1389 -143
rect 1409 -147 1411 -139
rect 1431 -147 1433 -143
rect 1447 -147 1449 -143
rect 1483 -147 1485 -143
rect 1505 -147 1507 -139
rect 1527 -147 1529 -143
rect 1543 -147 1545 -143
rect 1574 -147 1576 -143
<< ptransistor >>
rect -523 265 -521 273
rect -504 265 -502 273
rect -485 265 -483 273
rect -463 257 -461 273
rect -441 265 -439 273
rect -425 265 -423 273
rect -389 265 -387 273
rect -367 257 -365 273
rect -345 265 -343 273
rect -329 265 -327 273
rect -298 265 -296 273
rect -273 265 -271 273
rect -254 265 -252 273
rect -232 257 -230 273
rect -210 265 -208 273
rect -194 265 -192 273
rect -158 265 -156 273
rect -136 257 -134 273
rect -114 265 -112 273
rect -98 265 -96 273
rect -67 265 -65 273
rect 22 265 24 273
rect 41 265 43 273
rect 63 257 65 273
rect 85 265 87 273
rect 101 265 103 273
rect 137 265 139 273
rect 159 257 161 273
rect 181 265 183 273
rect 197 265 199 273
rect 228 265 230 273
rect 360 265 362 273
rect 379 265 381 273
rect 401 257 403 273
rect 423 265 425 273
rect 439 265 441 273
rect 475 265 477 273
rect 497 257 499 273
rect 519 265 521 273
rect 535 265 537 273
rect 566 265 568 273
rect 613 265 615 273
rect 632 265 634 273
rect 654 257 656 273
rect 676 265 678 273
rect 692 265 694 273
rect 728 265 730 273
rect 750 257 752 273
rect 772 265 774 273
rect 788 265 790 273
rect 819 265 821 273
rect 877 265 879 273
rect 896 265 898 273
rect 918 257 920 273
rect 940 265 942 273
rect 956 265 958 273
rect 992 265 994 273
rect 1014 257 1016 273
rect 1036 265 1038 273
rect 1052 265 1054 273
rect 1083 265 1085 273
rect 1161 265 1163 273
rect 1180 265 1182 273
rect 1202 257 1204 273
rect 1224 265 1226 273
rect 1240 265 1242 273
rect 1276 265 1278 273
rect 1298 257 1300 273
rect 1320 265 1322 273
rect 1336 265 1338 273
rect 1367 265 1369 273
rect 1413 265 1415 273
rect 1432 265 1434 273
rect 1454 257 1456 273
rect 1476 265 1478 273
rect 1492 265 1494 273
rect 1528 265 1530 273
rect 1550 257 1552 273
rect 1572 265 1574 273
rect 1588 265 1590 273
rect 1619 265 1621 273
rect 1672 265 1674 273
rect 1691 265 1693 273
rect 1713 257 1715 273
rect 1735 265 1737 273
rect 1751 265 1753 273
rect 1787 265 1789 273
rect 1809 257 1811 273
rect 1831 265 1833 273
rect 1847 265 1849 273
rect 1878 265 1880 273
rect 6 98 8 106
rect 22 98 24 106
rect 38 90 40 106
rect 46 90 48 106
rect 54 90 56 106
rect 62 90 64 106
rect 81 98 83 106
rect 89 98 91 106
rect 107 98 109 106
rect 135 98 137 106
rect 151 98 153 106
rect 167 90 169 106
rect 175 90 177 106
rect 183 90 185 106
rect 191 90 193 106
rect 210 98 212 106
rect 218 98 220 106
rect 236 98 238 106
rect 263 98 265 106
rect 271 98 273 106
rect 289 98 291 106
rect 321 98 323 106
rect 337 98 339 106
rect 353 90 355 106
rect 361 90 363 106
rect 369 90 371 106
rect 377 90 379 106
rect 396 98 398 106
rect 404 98 406 106
rect 422 98 424 106
rect 450 98 452 106
rect 466 98 468 106
rect 482 90 484 106
rect 490 90 492 106
rect 498 90 500 106
rect 506 90 508 106
rect 525 98 527 106
rect 533 98 535 106
rect 551 98 553 106
rect 578 98 580 106
rect 586 98 588 106
rect 604 98 606 106
rect 885 98 887 106
rect 901 98 903 106
rect 917 90 919 106
rect 925 90 927 106
rect 933 90 935 106
rect 941 90 943 106
rect 960 98 962 106
rect 968 98 970 106
rect 986 98 988 106
rect 1014 98 1016 106
rect 1030 98 1032 106
rect 1046 90 1048 106
rect 1054 90 1056 106
rect 1062 90 1064 106
rect 1070 90 1072 106
rect 1089 98 1091 106
rect 1097 98 1099 106
rect 1115 98 1117 106
rect 1142 98 1144 106
rect 1150 98 1152 106
rect 1168 98 1170 106
rect 1468 98 1470 106
rect 1484 98 1486 106
rect 1500 90 1502 106
rect 1508 90 1510 106
rect 1516 90 1518 106
rect 1524 90 1526 106
rect 1543 98 1545 106
rect 1551 98 1553 106
rect 1569 98 1571 106
rect 1597 98 1599 106
rect 1613 98 1615 106
rect 1629 90 1631 106
rect 1637 90 1639 106
rect 1645 90 1647 106
rect 1653 90 1655 106
rect 1672 98 1674 106
rect 1680 98 1682 106
rect 1698 98 1700 106
rect 1725 98 1727 106
rect 1733 98 1735 106
rect 1751 98 1753 106
rect 10 -108 12 -100
rect 29 -108 31 -100
rect 51 -116 53 -100
rect 73 -108 75 -100
rect 89 -108 91 -100
rect 125 -108 127 -100
rect 147 -116 149 -100
rect 169 -108 171 -100
rect 185 -108 187 -100
rect 216 -108 218 -100
rect 256 -108 258 -100
rect 275 -108 277 -100
rect 297 -116 299 -100
rect 319 -108 321 -100
rect 335 -108 337 -100
rect 371 -108 373 -100
rect 393 -116 395 -100
rect 415 -108 417 -100
rect 431 -108 433 -100
rect 462 -108 464 -100
rect 757 -108 759 -100
rect 776 -108 778 -100
rect 798 -116 800 -100
rect 820 -108 822 -100
rect 836 -108 838 -100
rect 872 -108 874 -100
rect 894 -116 896 -100
rect 916 -108 918 -100
rect 932 -108 934 -100
rect 963 -108 965 -100
rect 1069 -108 1071 -100
rect 1088 -108 1090 -100
rect 1110 -116 1112 -100
rect 1132 -108 1134 -100
rect 1148 -108 1150 -100
rect 1184 -108 1186 -100
rect 1206 -116 1208 -100
rect 1228 -108 1230 -100
rect 1244 -108 1246 -100
rect 1275 -108 1277 -100
rect 1368 -108 1370 -100
rect 1387 -108 1389 -100
rect 1409 -116 1411 -100
rect 1431 -108 1433 -100
rect 1447 -108 1449 -100
rect 1483 -108 1485 -100
rect 1505 -116 1507 -100
rect 1527 -108 1529 -100
rect 1543 -108 1545 -100
rect 1574 -108 1576 -100
<< polycontact >>
rect -486 303 -482 307
rect -330 303 -326 307
rect -255 303 -251 307
rect -99 303 -95 307
rect 40 303 44 307
rect 196 303 200 307
rect 378 303 382 307
rect 534 303 538 307
rect 631 303 635 307
rect 787 303 791 307
rect 895 303 899 307
rect 1051 303 1055 307
rect 1179 303 1183 307
rect 1335 303 1339 307
rect 1431 303 1435 307
rect 1587 303 1591 307
rect 1690 303 1694 307
rect 1846 303 1850 307
rect -426 294 -422 298
rect -390 294 -386 298
rect -195 294 -191 298
rect -159 294 -155 298
rect 100 294 104 298
rect 136 294 140 298
rect 438 294 442 298
rect 474 294 478 298
rect 691 294 695 298
rect 727 294 731 298
rect 955 294 959 298
rect 991 294 995 298
rect 1239 294 1243 298
rect 1275 294 1279 298
rect 1491 294 1495 298
rect 1527 294 1531 298
rect 1750 294 1754 298
rect 1786 294 1790 298
rect -527 245 -523 249
rect -508 245 -504 249
rect -467 245 -463 249
rect -445 245 -441 249
rect -371 245 -367 249
rect -349 245 -345 249
rect -302 245 -298 249
rect -277 245 -273 249
rect -236 245 -232 249
rect -214 245 -210 249
rect -140 245 -136 249
rect -118 245 -114 249
rect -71 245 -67 249
rect 18 245 22 249
rect 59 245 63 249
rect 81 245 85 249
rect 155 245 159 249
rect 177 245 181 249
rect 224 245 228 249
rect 356 245 360 249
rect 397 245 401 249
rect 419 245 423 249
rect 493 245 497 249
rect 515 245 519 249
rect 562 245 566 249
rect 609 245 613 249
rect 650 245 654 249
rect 672 245 676 249
rect 746 245 750 249
rect 768 245 772 249
rect 815 245 819 249
rect 873 245 877 249
rect 914 245 918 249
rect 936 245 940 249
rect 1010 245 1014 249
rect 1032 245 1036 249
rect 1079 245 1083 249
rect 1157 245 1161 249
rect 1198 245 1202 249
rect 1220 245 1224 249
rect 1294 245 1298 249
rect 1316 245 1320 249
rect 1363 245 1367 249
rect 1409 245 1413 249
rect 1450 245 1454 249
rect 1472 245 1476 249
rect 1546 245 1550 249
rect 1568 245 1572 249
rect 1615 245 1619 249
rect 1668 245 1672 249
rect 1709 245 1713 249
rect 1731 245 1735 249
rect 1805 245 1809 249
rect 1827 245 1831 249
rect 1874 245 1878 249
rect -486 189 -482 193
rect -330 189 -326 193
rect -255 189 -251 193
rect -99 189 -95 193
rect 40 189 44 193
rect 196 189 200 193
rect 378 189 382 193
rect 534 189 538 193
rect 631 189 635 193
rect 787 189 791 193
rect 895 189 899 193
rect 1051 189 1055 193
rect 1179 189 1183 193
rect 1335 189 1339 193
rect 1431 189 1435 193
rect 1587 189 1591 193
rect 1690 189 1694 193
rect 1846 189 1850 193
rect -426 180 -422 184
rect -390 180 -386 184
rect -195 180 -191 184
rect -159 180 -155 184
rect 100 180 104 184
rect 136 180 140 184
rect 438 180 442 184
rect 474 180 478 184
rect 691 180 695 184
rect 727 180 731 184
rect 955 180 959 184
rect 991 180 995 184
rect 1239 180 1243 184
rect 1275 180 1279 184
rect 1491 180 1495 184
rect 1527 180 1531 184
rect 1750 180 1754 184
rect 1786 180 1790 184
rect 336 149 340 153
rect 150 133 154 137
rect 21 126 25 130
rect 5 119 9 123
rect 37 119 41 123
rect 53 119 57 123
rect 80 118 84 122
rect 134 119 138 123
rect 166 119 170 123
rect 182 119 186 123
rect 209 118 213 122
rect 320 119 324 123
rect 900 145 904 149
rect 465 135 469 139
rect 352 119 356 123
rect 368 119 372 123
rect 395 118 399 122
rect 449 119 453 123
rect 481 119 485 123
rect 497 119 501 123
rect 524 118 528 122
rect 884 119 888 123
rect 1483 144 1487 148
rect 1029 135 1033 139
rect 916 119 920 123
rect 932 119 936 123
rect 959 118 963 122
rect 1013 119 1017 123
rect 1045 119 1049 123
rect 1061 119 1065 123
rect 1088 118 1092 122
rect 1467 119 1471 123
rect 1612 135 1616 139
rect 1499 119 1503 123
rect 1515 119 1519 123
rect 1542 118 1546 122
rect 1596 119 1600 123
rect 1628 119 1632 123
rect 1644 119 1648 123
rect 1671 118 1675 122
rect 2 87 6 91
rect 103 63 107 67
rect 131 86 135 90
rect 147 86 151 90
rect 232 63 236 67
rect 259 63 263 67
rect 285 89 289 93
rect 333 86 337 90
rect 418 63 422 67
rect 21 17 25 21
rect 45 17 49 21
rect 61 17 65 21
rect 88 18 92 22
rect 446 86 450 90
rect 547 63 551 67
rect 574 63 578 67
rect 600 89 604 93
rect 897 86 901 90
rect 982 63 986 67
rect 150 17 154 21
rect 174 17 178 21
rect 190 17 194 21
rect 217 18 221 22
rect 270 18 274 22
rect 336 17 340 21
rect 360 17 364 21
rect 376 17 380 21
rect 403 18 407 22
rect 1010 86 1014 90
rect 1111 63 1115 67
rect 1138 63 1142 67
rect 1164 89 1168 93
rect 1565 63 1569 67
rect 465 17 469 21
rect 489 17 493 21
rect 505 17 509 21
rect 532 18 536 22
rect 585 18 589 22
rect 900 17 904 21
rect 924 17 928 21
rect 940 17 944 21
rect 967 18 971 22
rect 1593 86 1597 90
rect 1694 63 1698 67
rect 1721 63 1725 67
rect 1747 89 1751 93
rect 1029 17 1033 21
rect 1053 17 1057 21
rect 1069 17 1073 21
rect 1096 18 1100 22
rect 1149 18 1153 22
rect 1483 17 1487 21
rect 1507 17 1511 21
rect 1523 17 1527 21
rect 1550 18 1554 22
rect 1612 17 1616 21
rect 1636 17 1640 21
rect 1652 17 1656 21
rect 1679 18 1683 22
rect 1732 18 1736 22
rect 9 -57 13 -53
rect 28 -70 32 -66
rect 184 -70 188 -66
rect 274 -70 278 -66
rect 430 -70 434 -66
rect 775 -70 779 -66
rect 931 -70 935 -66
rect 1087 -70 1091 -66
rect 1243 -70 1247 -66
rect 1386 -70 1390 -66
rect 1542 -70 1546 -66
rect 88 -79 92 -75
rect 124 -79 128 -75
rect 334 -79 338 -75
rect 370 -79 374 -75
rect 835 -79 839 -75
rect 871 -79 875 -75
rect 1147 -79 1151 -75
rect 1183 -79 1187 -75
rect 1446 -79 1450 -75
rect 1482 -79 1486 -75
rect 47 -128 51 -124
rect 69 -128 73 -124
rect 143 -128 147 -124
rect 165 -128 169 -124
rect 212 -128 216 -124
rect 252 -128 256 -124
rect 293 -128 297 -124
rect 315 -128 319 -124
rect 389 -128 393 -124
rect 411 -128 415 -124
rect 458 -128 462 -124
rect 753 -128 757 -124
rect 794 -128 798 -124
rect 816 -128 820 -124
rect 890 -128 894 -124
rect 912 -128 916 -124
rect 959 -128 963 -124
rect 1065 -128 1069 -124
rect 1106 -128 1110 -124
rect 1128 -128 1132 -124
rect 1202 -128 1206 -124
rect 1224 -128 1228 -124
rect 1271 -128 1275 -124
rect 1364 -128 1368 -124
rect 1405 -128 1409 -124
rect 1427 -128 1431 -124
rect 1501 -128 1505 -124
rect 1523 -128 1527 -124
rect 1570 -128 1574 -124
rect 28 -184 32 -180
rect 184 -184 188 -180
rect 274 -184 278 -180
rect 430 -184 434 -180
rect 775 -184 779 -180
rect 931 -184 935 -180
rect 1087 -184 1091 -180
rect 1243 -184 1247 -180
rect 1386 -184 1390 -180
rect 1542 -184 1546 -180
rect 88 -193 92 -189
rect 124 -193 128 -189
rect 334 -193 338 -189
rect 370 -193 374 -189
rect 835 -193 839 -189
rect 871 -193 875 -189
rect 1147 -193 1151 -189
rect 1183 -193 1187 -189
rect 1446 -193 1450 -189
rect 1482 -193 1486 -189
<< ndcontact >>
rect -528 226 -524 230
rect -520 226 -516 230
rect -509 226 -505 230
rect -501 226 -497 230
rect -490 226 -486 230
rect -482 226 -478 230
rect -468 226 -464 234
rect -460 226 -456 234
rect -446 226 -442 230
rect -438 226 -434 230
rect -430 226 -426 230
rect -422 226 -418 230
rect -394 226 -390 230
rect -386 226 -382 230
rect -372 226 -368 234
rect -364 226 -360 234
rect -350 226 -346 230
rect -342 226 -338 230
rect -334 226 -330 230
rect -326 226 -322 230
rect -303 226 -299 230
rect -295 226 -291 230
rect -278 226 -274 230
rect -270 226 -266 230
rect -259 226 -255 230
rect -251 226 -247 230
rect -237 226 -233 234
rect -229 226 -225 234
rect -215 226 -211 230
rect -207 226 -203 230
rect -199 226 -195 230
rect -191 226 -187 230
rect -163 226 -159 230
rect -155 226 -151 230
rect -141 226 -137 234
rect -133 226 -129 234
rect -119 226 -115 230
rect -111 226 -107 230
rect -103 226 -99 230
rect -95 226 -91 230
rect -72 226 -68 230
rect -64 226 -60 230
rect 17 226 21 230
rect 25 226 29 230
rect 36 226 40 230
rect 44 226 48 230
rect 58 226 62 234
rect 66 226 70 234
rect 80 226 84 230
rect 88 226 92 230
rect 96 226 100 230
rect 104 226 108 230
rect 132 226 136 230
rect 140 226 144 230
rect 154 226 158 234
rect 162 226 166 234
rect 176 226 180 230
rect 184 226 188 230
rect 192 226 196 230
rect 200 226 204 230
rect 223 226 227 230
rect 231 226 235 230
rect 355 226 359 230
rect 363 226 367 230
rect 374 226 378 230
rect 382 226 386 230
rect 396 226 400 234
rect 404 226 408 234
rect 418 226 422 230
rect 426 226 430 230
rect 434 226 438 230
rect 442 226 446 230
rect 470 226 474 230
rect 478 226 482 230
rect 492 226 496 234
rect 500 226 504 234
rect 514 226 518 230
rect 522 226 526 230
rect 530 226 534 230
rect 538 226 542 230
rect 561 226 565 230
rect 569 226 573 230
rect 608 226 612 230
rect 616 226 620 230
rect 627 226 631 230
rect 635 226 639 230
rect 649 226 653 234
rect 657 226 661 234
rect 671 226 675 230
rect 679 226 683 230
rect 687 226 691 230
rect 695 226 699 230
rect 723 226 727 230
rect 731 226 735 230
rect 745 226 749 234
rect 753 226 757 234
rect 767 226 771 230
rect 775 226 779 230
rect 783 226 787 230
rect 791 226 795 230
rect 814 226 818 230
rect 822 226 826 230
rect 872 226 876 230
rect 880 226 884 230
rect 891 226 895 230
rect 899 226 903 230
rect 913 226 917 234
rect 921 226 925 234
rect 935 226 939 230
rect 943 226 947 230
rect 951 226 955 230
rect 959 226 963 230
rect 987 226 991 230
rect 995 226 999 230
rect 1009 226 1013 234
rect 1017 226 1021 234
rect 1031 226 1035 230
rect 1039 226 1043 230
rect 1047 226 1051 230
rect 1055 226 1059 230
rect 1078 226 1082 230
rect 1086 226 1090 230
rect 1156 226 1160 230
rect 1164 226 1168 230
rect 1175 226 1179 230
rect 1183 226 1187 230
rect 1197 226 1201 234
rect 1205 226 1209 234
rect 1219 226 1223 230
rect 1227 226 1231 230
rect 1235 226 1239 230
rect 1243 226 1247 230
rect 1271 226 1275 230
rect 1279 226 1283 230
rect 1293 226 1297 234
rect 1301 226 1305 234
rect 1315 226 1319 230
rect 1323 226 1327 230
rect 1331 226 1335 230
rect 1339 226 1343 230
rect 1362 226 1366 230
rect 1370 226 1374 230
rect 1408 226 1412 230
rect 1416 226 1420 230
rect 1427 226 1431 230
rect 1435 226 1439 230
rect 1449 226 1453 234
rect 1457 226 1461 234
rect 1471 226 1475 230
rect 1479 226 1483 230
rect 1487 226 1491 230
rect 1495 226 1499 230
rect 1523 226 1527 230
rect 1531 226 1535 230
rect 1545 226 1549 234
rect 1553 226 1557 234
rect 1567 226 1571 230
rect 1575 226 1579 230
rect 1583 226 1587 230
rect 1591 226 1595 230
rect 1614 226 1618 230
rect 1622 226 1626 230
rect 1667 226 1671 230
rect 1675 226 1679 230
rect 1686 226 1690 230
rect 1694 226 1698 230
rect 1708 226 1712 234
rect 1716 226 1720 234
rect 1730 226 1734 230
rect 1738 226 1742 230
rect 1746 226 1750 230
rect 1754 226 1758 230
rect 1782 226 1786 230
rect 1790 226 1794 230
rect 1804 226 1808 234
rect 1812 226 1816 234
rect 1826 226 1830 230
rect 1834 226 1838 230
rect 1842 226 1846 230
rect 1850 226 1854 230
rect 1873 226 1877 230
rect 1881 226 1885 230
rect 1 34 5 38
rect 9 34 13 38
rect 17 34 21 38
rect 25 34 29 38
rect 33 34 37 42
rect 49 34 53 42
rect 65 34 69 42
rect 74 34 78 42
rect 94 34 98 42
rect 102 34 106 38
rect 110 34 114 38
rect 130 34 134 38
rect 138 34 142 38
rect 146 34 150 38
rect 154 34 158 38
rect 162 34 166 42
rect 178 34 182 42
rect 194 34 198 42
rect 203 34 207 42
rect 223 34 227 42
rect 231 34 235 38
rect 239 34 243 38
rect 257 35 261 43
rect 266 35 270 43
rect 274 35 278 43
rect 283 34 287 38
rect 293 34 297 38
rect 316 34 320 38
rect 324 34 328 38
rect 332 34 336 38
rect 340 34 344 38
rect 348 34 352 42
rect 364 34 368 42
rect 380 34 384 42
rect 389 34 393 42
rect 409 34 413 42
rect 417 34 421 38
rect 425 34 429 38
rect 445 34 449 38
rect 453 34 457 38
rect 461 34 465 38
rect 469 34 473 38
rect 477 34 481 42
rect 493 34 497 42
rect 509 34 513 42
rect 518 34 522 42
rect 538 34 542 42
rect 546 34 550 38
rect 554 34 558 38
rect 572 35 576 43
rect 581 35 585 43
rect 589 35 593 43
rect 598 34 602 38
rect 608 34 612 38
rect 880 34 884 38
rect 888 34 892 38
rect 896 34 900 38
rect 904 34 908 38
rect 912 34 916 42
rect 928 34 932 42
rect 944 34 948 42
rect 953 34 957 42
rect 973 34 977 42
rect 981 34 985 38
rect 989 34 993 38
rect 1009 34 1013 38
rect 1017 34 1021 38
rect 1025 34 1029 38
rect 1033 34 1037 38
rect 1041 34 1045 42
rect 1057 34 1061 42
rect 1073 34 1077 42
rect 1082 34 1086 42
rect 1102 34 1106 42
rect 1110 34 1114 38
rect 1118 34 1122 38
rect 1136 35 1140 43
rect 1145 35 1149 43
rect 1153 35 1157 43
rect 1162 34 1166 38
rect 1172 34 1176 38
rect 1463 34 1467 38
rect 1471 34 1475 38
rect 1479 34 1483 38
rect 1487 34 1491 38
rect 1495 34 1499 42
rect 1511 34 1515 42
rect 1527 34 1531 42
rect 1536 34 1540 42
rect 1556 34 1560 42
rect 1564 34 1568 38
rect 1572 34 1576 38
rect 1592 34 1596 38
rect 1600 34 1604 38
rect 1608 34 1612 38
rect 1616 34 1620 38
rect 1624 34 1628 42
rect 1640 34 1644 42
rect 1656 34 1660 42
rect 1665 34 1669 42
rect 1685 34 1689 42
rect 1693 34 1697 38
rect 1701 34 1705 38
rect 1719 35 1723 43
rect 1728 35 1732 43
rect 1736 35 1740 43
rect 1745 34 1749 38
rect 1755 34 1759 38
rect 5 -147 9 -143
rect 13 -147 17 -143
rect 24 -147 28 -143
rect 32 -147 36 -143
rect 46 -147 50 -139
rect 54 -147 58 -139
rect 68 -147 72 -143
rect 76 -147 80 -143
rect 84 -147 88 -143
rect 92 -147 96 -143
rect 120 -147 124 -143
rect 128 -147 132 -143
rect 142 -147 146 -139
rect 150 -147 154 -139
rect 164 -147 168 -143
rect 172 -147 176 -143
rect 180 -147 184 -143
rect 188 -147 192 -143
rect 211 -147 215 -143
rect 219 -147 223 -143
rect 251 -147 255 -143
rect 259 -147 263 -143
rect 270 -147 274 -143
rect 278 -147 282 -143
rect 292 -147 296 -139
rect 300 -147 304 -139
rect 314 -147 318 -143
rect 322 -147 326 -143
rect 330 -147 334 -143
rect 338 -147 342 -143
rect 366 -147 370 -143
rect 374 -147 378 -143
rect 388 -147 392 -139
rect 396 -147 400 -139
rect 410 -147 414 -143
rect 418 -147 422 -143
rect 426 -147 430 -143
rect 434 -147 438 -143
rect 457 -147 461 -143
rect 465 -147 469 -143
rect 752 -147 756 -143
rect 760 -147 764 -143
rect 771 -147 775 -143
rect 779 -147 783 -143
rect 793 -147 797 -139
rect 801 -147 805 -139
rect 815 -147 819 -143
rect 823 -147 827 -143
rect 831 -147 835 -143
rect 839 -147 843 -143
rect 867 -147 871 -143
rect 875 -147 879 -143
rect 889 -147 893 -139
rect 897 -147 901 -139
rect 911 -147 915 -143
rect 919 -147 923 -143
rect 927 -147 931 -143
rect 935 -147 939 -143
rect 958 -147 962 -143
rect 966 -147 970 -143
rect 1064 -147 1068 -143
rect 1072 -147 1076 -143
rect 1083 -147 1087 -143
rect 1091 -147 1095 -143
rect 1105 -147 1109 -139
rect 1113 -147 1117 -139
rect 1127 -147 1131 -143
rect 1135 -147 1139 -143
rect 1143 -147 1147 -143
rect 1151 -147 1155 -143
rect 1179 -147 1183 -143
rect 1187 -147 1191 -143
rect 1201 -147 1205 -139
rect 1209 -147 1213 -139
rect 1223 -147 1227 -143
rect 1231 -147 1235 -143
rect 1239 -147 1243 -143
rect 1247 -147 1251 -143
rect 1270 -147 1274 -143
rect 1278 -147 1282 -143
rect 1363 -147 1367 -143
rect 1371 -147 1375 -143
rect 1382 -147 1386 -143
rect 1390 -147 1394 -143
rect 1404 -147 1408 -139
rect 1412 -147 1416 -139
rect 1426 -147 1430 -143
rect 1434 -147 1438 -143
rect 1442 -147 1446 -143
rect 1450 -147 1454 -143
rect 1478 -147 1482 -143
rect 1486 -147 1490 -143
rect 1500 -147 1504 -139
rect 1508 -147 1512 -139
rect 1522 -147 1526 -143
rect 1530 -147 1534 -143
rect 1538 -147 1542 -143
rect 1546 -147 1550 -143
rect 1569 -147 1573 -143
rect 1577 -147 1581 -143
<< pdcontact >>
rect -528 265 -524 273
rect -520 265 -516 273
rect -509 265 -505 273
rect -501 265 -497 273
rect -490 265 -486 273
rect -482 265 -478 273
rect -468 257 -464 273
rect -460 257 -456 273
rect -446 265 -442 273
rect -438 265 -434 273
rect -430 265 -426 273
rect -422 265 -418 273
rect -394 265 -390 273
rect -386 265 -382 273
rect -372 257 -368 273
rect -364 257 -360 273
rect -350 265 -346 273
rect -342 265 -338 273
rect -334 265 -330 273
rect -326 265 -322 273
rect -303 265 -299 273
rect -295 265 -291 273
rect -278 265 -274 273
rect -270 265 -266 273
rect -259 265 -255 273
rect -251 265 -247 273
rect -237 257 -233 273
rect -229 257 -225 273
rect -215 265 -211 273
rect -207 265 -203 273
rect -199 265 -195 273
rect -191 265 -187 273
rect -163 265 -159 273
rect -155 265 -151 273
rect -141 257 -137 273
rect -133 257 -129 273
rect -119 265 -115 273
rect -111 265 -107 273
rect -103 265 -99 273
rect -95 265 -91 273
rect -72 265 -68 273
rect -64 265 -60 273
rect 17 265 21 273
rect 25 265 29 273
rect 36 265 40 273
rect 44 265 48 273
rect 58 257 62 273
rect 66 257 70 273
rect 80 265 84 273
rect 88 265 92 273
rect 96 265 100 273
rect 104 265 108 273
rect 132 265 136 273
rect 140 265 144 273
rect 154 257 158 273
rect 162 257 166 273
rect 176 265 180 273
rect 184 265 188 273
rect 192 265 196 273
rect 200 265 204 273
rect 223 265 227 273
rect 231 265 235 273
rect 355 265 359 273
rect 363 265 367 273
rect 374 265 378 273
rect 382 265 386 273
rect 396 257 400 273
rect 404 257 408 273
rect 418 265 422 273
rect 426 265 430 273
rect 434 265 438 273
rect 442 265 446 273
rect 470 265 474 273
rect 478 265 482 273
rect 492 257 496 273
rect 500 257 504 273
rect 514 265 518 273
rect 522 265 526 273
rect 530 265 534 273
rect 538 265 542 273
rect 561 265 565 273
rect 569 265 573 273
rect 608 265 612 273
rect 616 265 620 273
rect 627 265 631 273
rect 635 265 639 273
rect 649 257 653 273
rect 657 257 661 273
rect 671 265 675 273
rect 679 265 683 273
rect 687 265 691 273
rect 695 265 699 273
rect 723 265 727 273
rect 731 265 735 273
rect 745 257 749 273
rect 753 257 757 273
rect 767 265 771 273
rect 775 265 779 273
rect 783 265 787 273
rect 791 265 795 273
rect 814 265 818 273
rect 822 265 826 273
rect 872 265 876 273
rect 880 265 884 273
rect 891 265 895 273
rect 899 265 903 273
rect 913 257 917 273
rect 921 257 925 273
rect 935 265 939 273
rect 943 265 947 273
rect 951 265 955 273
rect 959 265 963 273
rect 987 265 991 273
rect 995 265 999 273
rect 1009 257 1013 273
rect 1017 257 1021 273
rect 1031 265 1035 273
rect 1039 265 1043 273
rect 1047 265 1051 273
rect 1055 265 1059 273
rect 1078 265 1082 273
rect 1086 265 1090 273
rect 1156 265 1160 273
rect 1164 265 1168 273
rect 1175 265 1179 273
rect 1183 265 1187 273
rect 1197 257 1201 273
rect 1205 257 1209 273
rect 1219 265 1223 273
rect 1227 265 1231 273
rect 1235 265 1239 273
rect 1243 265 1247 273
rect 1271 265 1275 273
rect 1279 265 1283 273
rect 1293 257 1297 273
rect 1301 257 1305 273
rect 1315 265 1319 273
rect 1323 265 1327 273
rect 1331 265 1335 273
rect 1339 265 1343 273
rect 1362 265 1366 273
rect 1370 265 1374 273
rect 1408 265 1412 273
rect 1416 265 1420 273
rect 1427 265 1431 273
rect 1435 265 1439 273
rect 1449 257 1453 273
rect 1457 257 1461 273
rect 1471 265 1475 273
rect 1479 265 1483 273
rect 1487 265 1491 273
rect 1495 265 1499 273
rect 1523 265 1527 273
rect 1531 265 1535 273
rect 1545 257 1549 273
rect 1553 257 1557 273
rect 1567 265 1571 273
rect 1575 265 1579 273
rect 1583 265 1587 273
rect 1591 265 1595 273
rect 1614 265 1618 273
rect 1622 265 1626 273
rect 1667 265 1671 273
rect 1675 265 1679 273
rect 1686 265 1690 273
rect 1694 265 1698 273
rect 1708 257 1712 273
rect 1716 257 1720 273
rect 1730 265 1734 273
rect 1738 265 1742 273
rect 1746 265 1750 273
rect 1754 265 1758 273
rect 1782 265 1786 273
rect 1790 265 1794 273
rect 1804 257 1808 273
rect 1812 257 1816 273
rect 1826 265 1830 273
rect 1834 265 1838 273
rect 1842 265 1846 273
rect 1850 265 1854 273
rect 1873 265 1877 273
rect 1881 265 1885 273
rect 1 98 5 106
rect 9 98 13 106
rect 17 98 21 106
rect 25 98 29 106
rect 33 90 37 106
rect 41 98 45 106
rect 49 90 53 106
rect 57 90 61 98
rect 65 90 69 106
rect 75 100 79 104
rect 84 100 88 104
rect 93 100 97 104
rect 102 98 106 106
rect 110 98 114 106
rect 130 98 134 106
rect 138 98 142 106
rect 146 98 150 106
rect 154 98 158 106
rect 162 90 166 106
rect 170 98 174 106
rect 178 90 182 106
rect 186 90 190 98
rect 194 90 198 106
rect 204 100 208 104
rect 213 100 217 104
rect 222 100 226 104
rect 231 98 235 106
rect 239 98 243 106
rect 257 98 261 106
rect 274 98 278 106
rect 283 98 287 106
rect 293 98 297 106
rect 316 98 320 106
rect 324 98 328 106
rect 332 98 336 106
rect 340 98 344 106
rect 348 90 352 106
rect 356 98 360 106
rect 364 90 368 106
rect 372 90 376 98
rect 380 90 384 106
rect 390 100 394 104
rect 399 100 403 104
rect 408 100 412 104
rect 417 98 421 106
rect 425 98 429 106
rect 445 98 449 106
rect 453 98 457 106
rect 461 98 465 106
rect 469 98 473 106
rect 477 90 481 106
rect 485 98 489 106
rect 493 90 497 106
rect 501 90 505 98
rect 509 90 513 106
rect 519 100 523 104
rect 528 100 532 104
rect 537 100 541 104
rect 546 98 550 106
rect 554 98 558 106
rect 572 98 576 106
rect 589 98 593 106
rect 598 98 602 106
rect 608 98 612 106
rect 880 98 884 106
rect 888 98 892 106
rect 896 98 900 106
rect 904 98 908 106
rect 912 90 916 106
rect 920 98 924 106
rect 928 90 932 106
rect 936 90 940 98
rect 944 90 948 106
rect 954 100 958 104
rect 963 100 967 104
rect 972 100 976 104
rect 981 98 985 106
rect 989 98 993 106
rect 1009 98 1013 106
rect 1017 98 1021 106
rect 1025 98 1029 106
rect 1033 98 1037 106
rect 1041 90 1045 106
rect 1049 98 1053 106
rect 1057 90 1061 106
rect 1065 90 1069 98
rect 1073 90 1077 106
rect 1083 100 1087 104
rect 1092 100 1096 104
rect 1101 100 1105 104
rect 1110 98 1114 106
rect 1118 98 1122 106
rect 1136 98 1140 106
rect 1153 98 1157 106
rect 1162 98 1166 106
rect 1172 98 1176 106
rect 1463 98 1467 106
rect 1471 98 1475 106
rect 1479 98 1483 106
rect 1487 98 1491 106
rect 1495 90 1499 106
rect 1503 98 1507 106
rect 1511 90 1515 106
rect 1519 90 1523 98
rect 1527 90 1531 106
rect 1537 100 1541 104
rect 1546 100 1550 104
rect 1555 100 1559 104
rect 1564 98 1568 106
rect 1572 98 1576 106
rect 1592 98 1596 106
rect 1600 98 1604 106
rect 1608 98 1612 106
rect 1616 98 1620 106
rect 1624 90 1628 106
rect 1632 98 1636 106
rect 1640 90 1644 106
rect 1648 90 1652 98
rect 1656 90 1660 106
rect 1666 100 1670 104
rect 1675 100 1679 104
rect 1684 100 1688 104
rect 1693 98 1697 106
rect 1701 98 1705 106
rect 1719 98 1723 106
rect 1736 98 1740 106
rect 1745 98 1749 106
rect 1755 98 1759 106
rect 5 -108 9 -100
rect 13 -108 17 -100
rect 24 -108 28 -100
rect 32 -108 36 -100
rect 46 -116 50 -100
rect 54 -116 58 -100
rect 68 -108 72 -100
rect 76 -108 80 -100
rect 84 -108 88 -100
rect 92 -108 96 -100
rect 120 -108 124 -100
rect 128 -108 132 -100
rect 142 -116 146 -100
rect 150 -116 154 -100
rect 164 -108 168 -100
rect 172 -108 176 -100
rect 180 -108 184 -100
rect 188 -108 192 -100
rect 211 -108 215 -100
rect 219 -108 223 -100
rect 251 -108 255 -100
rect 259 -108 263 -100
rect 270 -108 274 -100
rect 278 -108 282 -100
rect 292 -116 296 -100
rect 300 -116 304 -100
rect 314 -108 318 -100
rect 322 -108 326 -100
rect 330 -108 334 -100
rect 338 -108 342 -100
rect 366 -108 370 -100
rect 374 -108 378 -100
rect 388 -116 392 -100
rect 396 -116 400 -100
rect 410 -108 414 -100
rect 418 -108 422 -100
rect 426 -108 430 -100
rect 434 -108 438 -100
rect 457 -108 461 -100
rect 465 -108 469 -100
rect 752 -108 756 -100
rect 760 -108 764 -100
rect 771 -108 775 -100
rect 779 -108 783 -100
rect 793 -116 797 -100
rect 801 -116 805 -100
rect 815 -108 819 -100
rect 823 -108 827 -100
rect 831 -108 835 -100
rect 839 -108 843 -100
rect 867 -108 871 -100
rect 875 -108 879 -100
rect 889 -116 893 -100
rect 897 -116 901 -100
rect 911 -108 915 -100
rect 919 -108 923 -100
rect 927 -108 931 -100
rect 935 -108 939 -100
rect 958 -108 962 -100
rect 966 -108 970 -100
rect 1064 -108 1068 -100
rect 1072 -108 1076 -100
rect 1083 -108 1087 -100
rect 1091 -108 1095 -100
rect 1105 -116 1109 -100
rect 1113 -116 1117 -100
rect 1127 -108 1131 -100
rect 1135 -108 1139 -100
rect 1143 -108 1147 -100
rect 1151 -108 1155 -100
rect 1179 -108 1183 -100
rect 1187 -108 1191 -100
rect 1201 -116 1205 -100
rect 1209 -116 1213 -100
rect 1223 -108 1227 -100
rect 1231 -108 1235 -100
rect 1239 -108 1243 -100
rect 1247 -108 1251 -100
rect 1270 -108 1274 -100
rect 1278 -108 1282 -100
rect 1363 -108 1367 -100
rect 1371 -108 1375 -100
rect 1382 -108 1386 -100
rect 1390 -108 1394 -100
rect 1404 -116 1408 -100
rect 1412 -116 1416 -100
rect 1426 -108 1430 -100
rect 1434 -108 1438 -100
rect 1442 -108 1446 -100
rect 1450 -108 1454 -100
rect 1478 -108 1482 -100
rect 1486 -108 1490 -100
rect 1500 -116 1504 -100
rect 1508 -116 1512 -100
rect 1522 -108 1526 -100
rect 1530 -108 1534 -100
rect 1538 -108 1542 -100
rect 1546 -108 1550 -100
rect 1569 -108 1573 -100
rect 1577 -108 1581 -100
<< m2contact >>
rect -519 293 -514 298
rect 1952 274 1960 282
rect -520 245 -515 250
rect -482 245 -477 250
rect -453 245 -449 249
rect -422 245 -417 250
rect -395 245 -390 250
rect -378 245 -373 250
rect -357 245 -352 250
rect -326 245 -321 250
rect -312 245 -307 250
rect -287 244 -282 249
rect -251 245 -246 250
rect -222 245 -218 249
rect -191 245 -186 250
rect -164 245 -159 250
rect -147 245 -142 250
rect -126 245 -121 250
rect -95 245 -90 250
rect -81 245 -76 250
rect -53 245 -48 250
rect 44 245 49 250
rect 73 245 77 249
rect 104 245 109 250
rect 131 245 136 250
rect 148 245 153 250
rect 169 245 174 250
rect 200 245 205 250
rect 214 245 219 250
rect 239 245 244 250
rect 382 245 387 250
rect 411 245 415 249
rect 442 245 447 250
rect 469 245 474 250
rect 486 245 491 250
rect 507 245 512 250
rect 538 245 543 250
rect 552 245 557 250
rect 577 245 582 250
rect 635 245 640 250
rect 664 245 668 249
rect 695 245 700 250
rect 722 245 727 250
rect 739 245 744 250
rect 760 245 765 250
rect 791 245 796 250
rect 805 245 810 250
rect 834 245 839 250
rect 899 245 904 250
rect 928 245 932 249
rect 959 245 964 250
rect 986 245 991 250
rect 1003 245 1008 250
rect 1024 245 1029 250
rect 1055 245 1060 250
rect 1069 245 1074 250
rect 1104 245 1109 250
rect 1183 245 1188 250
rect 1212 245 1216 249
rect 1243 245 1248 250
rect 1270 245 1275 250
rect 1287 245 1292 250
rect 1308 245 1313 250
rect 1339 245 1344 250
rect 1353 245 1358 250
rect 1384 245 1389 250
rect 1435 245 1440 250
rect 1464 245 1468 249
rect 1495 245 1500 250
rect 1522 245 1527 250
rect 1539 245 1544 250
rect 1560 245 1565 250
rect 1591 245 1596 250
rect 1605 245 1610 250
rect 1636 245 1641 250
rect 1694 245 1699 250
rect 1723 245 1727 249
rect 1754 245 1759 250
rect 1781 245 1786 250
rect 1798 245 1803 250
rect 1819 245 1824 250
rect 1850 245 1855 250
rect 1864 245 1869 250
rect 1891 245 1896 250
rect -519 189 -514 194
rect 320 160 325 165
rect 1467 160 1472 165
rect 149 141 154 146
rect 20 133 25 138
rect 45 119 50 124
rect 174 119 179 124
rect 349 148 354 153
rect 883 151 888 156
rect 458 135 463 140
rect 360 119 365 124
rect 489 119 494 124
rect 900 152 905 157
rect 1021 134 1026 139
rect 924 119 929 124
rect 1053 119 1058 124
rect 1482 150 1487 155
rect 1605 135 1610 140
rect 1507 119 1512 124
rect 1636 119 1641 124
rect 1770 109 1778 117
rect -6 87 -1 92
rect 9 65 14 70
rect 25 65 30 70
rect 69 71 74 76
rect 124 85 129 90
rect 117 62 122 67
rect 138 65 143 70
rect 154 65 159 70
rect 198 71 203 76
rect 301 89 306 94
rect 324 65 329 70
rect 340 65 345 70
rect 384 71 389 76
rect 439 85 444 90
rect 432 62 437 67
rect 453 65 458 70
rect 469 65 474 70
rect 513 71 518 76
rect 616 89 621 94
rect 888 65 893 70
rect 904 65 909 70
rect 948 71 953 76
rect 1003 85 1008 90
rect 996 62 1001 67
rect 1017 65 1022 70
rect 1033 65 1038 70
rect 1077 71 1082 76
rect 1180 89 1185 94
rect 1471 65 1476 70
rect 1487 65 1492 70
rect 1531 71 1536 76
rect 1586 85 1591 90
rect 1579 62 1584 67
rect 1600 65 1605 70
rect 1616 65 1621 70
rect 1660 71 1665 76
rect 1802 54 1807 59
rect 53 16 58 21
rect 182 16 187 21
rect 269 11 274 16
rect 368 16 373 21
rect 497 16 502 21
rect 584 11 589 16
rect 932 16 937 21
rect 1061 16 1066 21
rect 1148 11 1153 16
rect 1515 16 1520 21
rect 1644 16 1649 21
rect 1731 11 1736 16
rect 1802 -3 1807 2
rect 1339 -40 1344 -35
rect 9 -49 14 -44
rect -9 -80 -4 -75
rect 1581 -97 1589 -89
rect 32 -128 37 -123
rect 61 -128 65 -124
rect 92 -128 97 -123
rect 119 -128 124 -123
rect 136 -128 141 -123
rect 157 -128 162 -123
rect 188 -128 193 -123
rect 202 -128 207 -123
rect 245 -128 250 -123
rect 278 -128 283 -123
rect 307 -128 311 -124
rect 338 -128 343 -123
rect 365 -128 370 -123
rect 382 -128 387 -123
rect 403 -128 408 -123
rect 434 -128 439 -123
rect 448 -128 453 -123
rect 739 -128 744 -123
rect 779 -128 784 -123
rect 808 -128 812 -124
rect 839 -128 844 -123
rect 866 -128 871 -123
rect 883 -128 888 -123
rect 904 -128 909 -123
rect 935 -128 940 -123
rect 949 -128 954 -123
rect 1042 -128 1047 -123
rect 1091 -128 1096 -123
rect 1120 -128 1124 -124
rect 1151 -128 1156 -123
rect 1178 -128 1183 -123
rect 1195 -128 1200 -123
rect 1216 -128 1221 -123
rect 1247 -128 1252 -123
rect 1261 -128 1266 -123
rect 1339 -128 1344 -123
rect 1390 -128 1395 -123
rect 1419 -128 1423 -124
rect 1450 -128 1455 -123
rect 1477 -128 1482 -123
rect 1494 -128 1499 -123
rect 1515 -128 1520 -123
rect 1546 -128 1551 -123
rect 1560 -128 1565 -123
rect -2 -184 3 -179
<< psubstratepcontact >>
rect -527 218 -523 222
rect -508 218 -504 222
rect -467 218 -463 222
rect -445 218 -441 222
rect -371 218 -367 222
rect -349 218 -345 222
rect -302 218 -298 222
rect -277 218 -273 222
rect -236 218 -232 222
rect -214 218 -210 222
rect -140 218 -136 222
rect -118 218 -114 222
rect -71 218 -67 222
rect 18 218 22 222
rect 59 218 63 222
rect 81 218 85 222
rect 155 218 159 222
rect 177 218 181 222
rect 224 218 228 222
rect 356 218 360 222
rect 397 218 401 222
rect 419 218 423 222
rect 493 218 497 222
rect 515 218 519 222
rect 562 218 566 222
rect 609 218 613 222
rect 650 218 654 222
rect 672 218 676 222
rect 746 218 750 222
rect 768 218 772 222
rect 815 218 819 222
rect 873 218 877 222
rect 914 218 918 222
rect 936 218 940 222
rect 1010 218 1014 222
rect 1032 218 1036 222
rect 1079 218 1083 222
rect 1157 218 1161 222
rect 1198 218 1202 222
rect 1220 218 1224 222
rect 1294 218 1298 222
rect 1316 218 1320 222
rect 1363 218 1367 222
rect 1409 218 1413 222
rect 1450 218 1454 222
rect 1472 218 1476 222
rect 1546 218 1550 222
rect 1568 218 1572 222
rect 1615 218 1619 222
rect 1668 218 1672 222
rect 1709 218 1713 222
rect 1731 218 1735 222
rect 1805 218 1809 222
rect 1827 218 1831 222
rect 1874 218 1878 222
rect 2 26 6 30
rect 75 26 79 30
rect 93 26 97 30
rect 103 26 107 30
rect 131 26 135 30
rect 204 26 208 30
rect 222 26 226 30
rect 232 26 236 30
rect 265 26 269 30
rect 283 26 287 30
rect 317 26 321 30
rect 390 26 394 30
rect 408 26 412 30
rect 418 26 422 30
rect 446 26 450 30
rect 519 26 523 30
rect 537 26 541 30
rect 547 26 551 30
rect 580 26 584 30
rect 598 26 602 30
rect 881 26 885 30
rect 954 26 958 30
rect 972 26 976 30
rect 982 26 986 30
rect 1010 26 1014 30
rect 1083 26 1087 30
rect 1101 26 1105 30
rect 1111 26 1115 30
rect 1144 26 1148 30
rect 1162 26 1166 30
rect 1464 26 1468 30
rect 1537 26 1541 30
rect 1555 26 1559 30
rect 1565 26 1569 30
rect 1593 26 1597 30
rect 1666 26 1670 30
rect 1684 26 1688 30
rect 1694 26 1698 30
rect 1727 26 1731 30
rect 1745 26 1749 30
rect 6 -155 10 -151
rect 47 -155 51 -151
rect 69 -155 73 -151
rect 143 -155 147 -151
rect 165 -155 169 -151
rect 212 -155 216 -151
rect 252 -155 256 -151
rect 293 -155 297 -151
rect 315 -155 319 -151
rect 389 -155 393 -151
rect 411 -155 415 -151
rect 458 -155 462 -151
rect 753 -155 757 -151
rect 794 -155 798 -151
rect 816 -155 820 -151
rect 890 -155 894 -151
rect 912 -155 916 -151
rect 959 -155 963 -151
rect 1065 -155 1069 -151
rect 1106 -155 1110 -151
rect 1128 -155 1132 -151
rect 1202 -155 1206 -151
rect 1224 -155 1228 -151
rect 1271 -155 1275 -151
rect 1364 -155 1368 -151
rect 1405 -155 1409 -151
rect 1427 -155 1431 -151
rect 1501 -155 1505 -151
rect 1523 -155 1527 -151
rect 1570 -155 1574 -151
<< nsubstratencontact >>
rect -527 277 -523 281
rect -508 277 -504 281
rect -467 277 -463 281
rect -445 277 -441 281
rect -371 277 -367 281
rect -349 277 -345 281
rect -302 277 -298 281
rect -277 277 -273 281
rect -236 277 -232 281
rect -214 277 -210 281
rect -140 277 -136 281
rect -118 277 -114 281
rect -71 277 -67 281
rect 18 277 22 281
rect 59 277 63 281
rect 81 277 85 281
rect 155 277 159 281
rect 177 277 181 281
rect 224 277 228 281
rect 356 277 360 281
rect 397 277 401 281
rect 419 277 423 281
rect 493 277 497 281
rect 515 277 519 281
rect 562 277 566 281
rect 609 277 613 281
rect 650 277 654 281
rect 672 277 676 281
rect 746 277 750 281
rect 768 277 772 281
rect 815 277 819 281
rect 873 277 877 281
rect 914 277 918 281
rect 936 277 940 281
rect 1010 277 1014 281
rect 1032 277 1036 281
rect 1079 277 1083 281
rect 1157 277 1161 281
rect 1198 277 1202 281
rect 1220 277 1224 281
rect 1294 277 1298 281
rect 1316 277 1320 281
rect 1363 277 1367 281
rect 1409 277 1413 281
rect 1450 277 1454 281
rect 1472 277 1476 281
rect 1546 277 1550 281
rect 1568 277 1572 281
rect 1615 277 1619 281
rect 1668 277 1672 281
rect 1709 277 1713 281
rect 1731 277 1735 281
rect 1805 277 1809 281
rect 1827 277 1831 281
rect 1874 277 1878 281
rect 15 110 19 114
rect 76 110 80 114
rect 93 110 97 114
rect 143 110 147 114
rect 205 110 209 114
rect 222 110 226 114
rect 258 110 262 114
rect 283 110 287 114
rect 330 110 334 114
rect 391 110 395 114
rect 408 110 412 114
rect 460 110 464 114
rect 520 110 524 114
rect 537 110 541 114
rect 573 110 577 114
rect 598 110 602 114
rect 895 110 899 114
rect 955 110 959 114
rect 972 110 976 114
rect 1024 110 1028 114
rect 1084 110 1088 114
rect 1101 110 1105 114
rect 1137 110 1141 114
rect 1162 110 1166 114
rect 1477 110 1481 114
rect 1538 110 1542 114
rect 1555 110 1559 114
rect 1607 110 1611 114
rect 1667 110 1671 114
rect 1684 110 1688 114
rect 1720 110 1724 114
rect 1745 110 1749 114
rect 4 -96 8 -92
rect 47 -96 51 -92
rect 69 -96 73 -92
rect 143 -96 147 -92
rect 165 -96 169 -92
rect 212 -96 216 -92
rect 252 -96 256 -92
rect 293 -96 297 -92
rect 315 -96 319 -92
rect 389 -96 393 -92
rect 411 -96 415 -92
rect 458 -96 462 -92
rect 753 -96 757 -92
rect 794 -96 798 -92
rect 816 -96 820 -92
rect 890 -96 894 -92
rect 912 -96 916 -92
rect 959 -96 963 -92
rect 1065 -96 1069 -92
rect 1106 -96 1110 -92
rect 1128 -96 1132 -92
rect 1202 -96 1206 -92
rect 1224 -96 1228 -92
rect 1271 -96 1275 -92
rect 1364 -96 1368 -92
rect 1405 -96 1409 -92
rect 1427 -96 1431 -92
rect 1501 -96 1505 -92
rect 1523 -96 1527 -92
rect 1570 -96 1574 -92
<< labels >>
rlabel polycontact -525 246 -525 246 1 clk
rlabel m2contact -517 248 -517 248 1 clkbar
rlabel polycontact -506 247 -506 247 1 A1
rlabel polycontact -276 247 -276 247 1 B1
rlabel polycontact 20 247 20 247 1 Cin
rlabel polycontact 4 89 4 89 1 A1bar
rlabel polycontact 22 128 22 128 1 B1bar
rlabel polycontact 152 135 152 135 1 Cinbar
rlabel polycontact 357 247 357 247 1 A2
rlabel polycontact 611 247 611 247 1 B2
rlabel polycontact 322 121 322 121 1 A2bar
rlabel polycontact 338 151 338 151 1 B2bar
rlabel polycontact 875 247 875 247 1 A3
rlabel polycontact 886 121 886 121 1 A3bar
rlabel polycontact 902 147 902 147 1 B3bar
rlabel polycontact 1159 247 1159 247 1 B3
rlabel polycontact 1411 247 1411 247 1 A4
rlabel polycontact 1670 247 1670 247 1 B4
rlabel polycontact 1469 121 1469 121 1 A4bar
rlabel polycontact 1485 145 1485 145 1 B4bar
rlabel polycontact 11 -55 11 -55 1 S0bar
rlabel metal1 225 -126 225 -126 1 S0
rlabel polycontact 254 -126 254 -126 1 S1bar
rlabel metal1 471 -126 471 -126 1 S1
rlabel polycontact 755 -126 755 -126 1 S2bar
rlabel metal1 972 -126 972 -126 1 S2
rlabel polycontact 1067 -126 1067 -126 1 S3bar
rlabel metal1 1284 -126 1284 -126 1 S3
rlabel polycontact 1366 -126 1366 -126 1 S4bar
rlabel metal1 1583 -126 1583 -126 1 S4
rlabel metal1 788 111 788 111 1 VDD
rlabel metal1 779 27 779 27 1 GND
<< end >>
