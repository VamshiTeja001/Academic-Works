magic
tech scmos
timestamp 1701919502
<< polysilicon >>
rect -46 35 -44 47
rect -28 35 -26 54
rect -10 35 -8 47
rect -2 35 0 37
rect 6 35 8 47
rect 14 35 16 37
rect 35 35 37 77
rect 53 35 55 84
rect 71 35 73 47
rect 79 35 81 37
rect 87 35 89 47
rect 95 35 97 37
rect 117 35 119 55
rect 125 35 127 55
rect 141 35 143 37
rect 168 35 170 77
rect 176 35 178 84
rect 192 35 194 37
rect 214 35 216 47
rect 222 35 224 37
rect 238 35 240 37
rect 262 35 264 47
rect 280 35 282 54
rect 298 35 300 47
rect 306 35 308 37
rect 314 35 316 47
rect 322 35 324 37
rect 343 35 345 77
rect 361 35 363 84
rect 379 35 381 47
rect 387 35 389 37
rect 395 35 397 47
rect 403 35 405 37
rect 425 35 427 55
rect 433 35 435 55
rect 449 35 451 37
rect 476 35 478 77
rect 484 35 486 84
rect 500 35 502 37
rect 522 35 524 47
rect 530 35 532 37
rect 546 35 548 37
rect 571 35 573 47
rect 589 35 591 54
rect 607 35 609 47
rect 615 35 617 37
rect 623 35 625 47
rect 631 35 633 37
rect 652 35 654 77
rect 670 35 672 84
rect 688 35 690 47
rect 696 35 698 37
rect 704 35 706 47
rect 712 35 714 37
rect 734 35 736 55
rect 742 35 744 55
rect 758 35 760 37
rect 785 35 787 77
rect 793 35 795 84
rect 809 35 811 37
rect 831 35 833 47
rect 839 35 841 37
rect 855 35 857 37
rect 890 35 892 47
rect 908 35 910 54
rect 926 35 928 47
rect 934 35 936 37
rect 942 35 944 47
rect 950 35 952 37
rect 971 35 973 77
rect 989 35 991 84
rect 1007 35 1009 47
rect 1015 35 1017 37
rect 1023 35 1025 47
rect 1031 35 1033 37
rect 1053 35 1055 55
rect 1061 35 1063 55
rect 1077 35 1079 37
rect 1104 35 1106 77
rect 1112 35 1114 84
rect 1128 35 1130 37
rect 1150 35 1152 47
rect 1158 35 1160 37
rect 1174 35 1176 37
rect 1198 35 1200 37
rect 1222 35 1224 37
rect 1248 35 1250 37
rect 1273 35 1275 37
rect -46 -15 -44 27
rect -28 -15 -26 27
rect -10 -11 -8 19
rect -2 -11 0 19
rect 6 -11 8 19
rect 14 -11 16 19
rect 35 -15 37 27
rect 53 -15 55 27
rect 71 -11 73 19
rect 79 -11 81 19
rect 87 -11 89 19
rect 95 -11 97 19
rect 117 -11 119 27
rect 125 -11 127 27
rect 141 -15 143 27
rect 168 -11 170 27
rect 176 -11 178 27
rect 192 -15 194 27
rect 214 -11 216 27
rect 222 -11 224 27
rect 238 -15 240 27
rect 262 -15 264 27
rect 280 -15 282 27
rect 298 -11 300 19
rect 306 -11 308 19
rect 314 -11 316 19
rect 322 -11 324 19
rect 343 -15 345 27
rect 361 -15 363 27
rect 379 -11 381 19
rect 387 -11 389 19
rect 395 -11 397 19
rect 403 -11 405 19
rect 425 -11 427 27
rect 433 -11 435 27
rect 449 -15 451 27
rect 476 -11 478 27
rect 484 -11 486 27
rect 500 -15 502 27
rect 522 -11 524 27
rect 530 -11 532 27
rect 546 -15 548 27
rect 571 -15 573 27
rect 589 -15 591 27
rect 607 -11 609 19
rect 615 -11 617 19
rect 623 -11 625 19
rect 631 -11 633 19
rect 652 -15 654 27
rect 670 -15 672 27
rect 688 -11 690 19
rect 696 -11 698 19
rect 704 -11 706 19
rect 712 -11 714 19
rect 734 -11 736 27
rect 742 -11 744 27
rect 758 -15 760 27
rect 785 -11 787 27
rect 793 -11 795 27
rect 809 -15 811 27
rect 831 -11 833 27
rect 839 -11 841 27
rect 855 -15 857 27
rect 890 -15 892 27
rect 908 -15 910 27
rect 926 -11 928 19
rect 934 -11 936 19
rect 942 -11 944 19
rect 950 -11 952 19
rect 971 -15 973 27
rect 989 -15 991 27
rect 1007 -11 1009 19
rect 1015 -11 1017 19
rect 1023 -11 1025 19
rect 1031 -11 1033 19
rect 1053 -11 1055 27
rect 1061 -11 1063 27
rect 1077 -15 1079 27
rect 1104 -11 1106 27
rect 1112 -11 1114 27
rect 1128 -15 1130 27
rect 1150 -11 1152 27
rect 1158 -11 1160 27
rect 1174 -15 1176 27
rect 1198 -15 1200 27
rect 1222 -15 1224 27
rect 1248 -15 1250 27
rect 1273 -15 1275 27
rect -46 -21 -44 -19
rect -28 -31 -26 -19
rect -10 -21 -8 -19
rect -2 -31 0 -19
rect 6 -21 8 -19
rect 14 -31 16 -19
rect 35 -21 37 -19
rect 53 -31 55 -19
rect 71 -21 73 -19
rect 79 -31 81 -19
rect 87 -21 89 -19
rect 95 -31 97 -19
rect 117 -21 119 -19
rect 125 -21 127 -19
rect 141 -21 143 -19
rect 168 -21 170 -19
rect 176 -21 178 -19
rect 192 -21 194 -19
rect 214 -21 216 -19
rect 222 -31 224 -19
rect 238 -21 240 -19
rect 262 -21 264 -19
rect 280 -31 282 -19
rect 298 -21 300 -19
rect 306 -31 308 -19
rect 314 -21 316 -19
rect 322 -31 324 -19
rect 343 -21 345 -19
rect 361 -31 363 -19
rect 379 -21 381 -19
rect 387 -31 389 -19
rect 395 -21 397 -19
rect 403 -31 405 -19
rect 425 -21 427 -19
rect 433 -21 435 -19
rect 449 -21 451 -19
rect 476 -21 478 -19
rect 484 -21 486 -19
rect 500 -21 502 -19
rect 522 -21 524 -19
rect 530 -31 532 -19
rect 546 -21 548 -19
rect 571 -21 573 -19
rect 589 -31 591 -19
rect 607 -21 609 -19
rect 615 -31 617 -19
rect 623 -21 625 -19
rect 631 -31 633 -19
rect 652 -21 654 -19
rect 670 -31 672 -19
rect 688 -21 690 -19
rect 696 -31 698 -19
rect 704 -21 706 -19
rect 712 -31 714 -19
rect 734 -21 736 -19
rect 742 -21 744 -19
rect 758 -21 760 -19
rect 785 -21 787 -19
rect 793 -21 795 -19
rect 809 -21 811 -19
rect 831 -21 833 -19
rect 839 -31 841 -19
rect 855 -21 857 -19
rect 890 -21 892 -19
rect 908 -31 910 -19
rect 926 -21 928 -19
rect 934 -31 936 -19
rect 942 -21 944 -19
rect 950 -31 952 -19
rect 971 -21 973 -19
rect 989 -31 991 -19
rect 1007 -21 1009 -19
rect 1015 -31 1017 -19
rect 1023 -21 1025 -19
rect 1031 -31 1033 -19
rect 1053 -21 1055 -19
rect 1061 -21 1063 -19
rect 1077 -21 1079 -19
rect 1104 -21 1106 -19
rect 1112 -21 1114 -19
rect 1128 -21 1130 -19
rect 1150 -21 1152 -19
rect 1158 -31 1160 -19
rect 1174 -21 1176 -19
rect 1198 -21 1200 -19
rect 1222 -21 1224 -19
rect 1248 -21 1250 -19
rect 1273 -21 1275 -19
<< ndiffusion >>
rect -47 -19 -46 -15
rect -44 -19 -43 -15
rect -29 -19 -28 -15
rect -26 -19 -25 -15
rect -11 -19 -10 -11
rect -8 -19 -2 -11
rect 0 -19 1 -11
rect 5 -19 6 -11
rect 8 -19 14 -11
rect 16 -19 17 -11
rect 34 -19 35 -15
rect 37 -19 38 -15
rect 52 -19 53 -15
rect 55 -19 56 -15
rect 70 -19 71 -11
rect 73 -19 79 -11
rect 81 -19 82 -11
rect 86 -19 87 -11
rect 89 -19 95 -11
rect 97 -19 98 -11
rect 116 -19 117 -11
rect 119 -19 125 -11
rect 127 -19 128 -11
rect 140 -19 141 -15
rect 143 -19 144 -15
rect 167 -19 168 -11
rect 170 -19 176 -11
rect 178 -19 179 -11
rect 191 -19 192 -15
rect 194 -19 195 -15
rect 213 -19 214 -11
rect 216 -19 217 -11
rect 221 -19 222 -11
rect 224 -19 225 -11
rect 237 -19 238 -15
rect 240 -19 241 -15
rect 261 -19 262 -15
rect 264 -19 265 -15
rect 279 -19 280 -15
rect 282 -19 283 -15
rect 297 -19 298 -11
rect 300 -19 306 -11
rect 308 -19 309 -11
rect 313 -19 314 -11
rect 316 -19 322 -11
rect 324 -19 325 -11
rect 342 -19 343 -15
rect 345 -19 346 -15
rect 360 -19 361 -15
rect 363 -19 364 -15
rect 378 -19 379 -11
rect 381 -19 387 -11
rect 389 -19 390 -11
rect 394 -19 395 -11
rect 397 -19 403 -11
rect 405 -19 406 -11
rect 424 -19 425 -11
rect 427 -19 433 -11
rect 435 -19 436 -11
rect 448 -19 449 -15
rect 451 -19 452 -15
rect 475 -19 476 -11
rect 478 -19 484 -11
rect 486 -19 487 -11
rect 499 -19 500 -15
rect 502 -19 503 -15
rect 521 -19 522 -11
rect 524 -19 525 -11
rect 529 -19 530 -11
rect 532 -19 533 -11
rect 545 -19 546 -15
rect 548 -19 549 -15
rect 570 -19 571 -15
rect 573 -19 574 -15
rect 588 -19 589 -15
rect 591 -19 592 -15
rect 606 -19 607 -11
rect 609 -19 615 -11
rect 617 -19 618 -11
rect 622 -19 623 -11
rect 625 -19 631 -11
rect 633 -19 634 -11
rect 651 -19 652 -15
rect 654 -19 655 -15
rect 669 -19 670 -15
rect 672 -19 673 -15
rect 687 -19 688 -11
rect 690 -19 696 -11
rect 698 -19 699 -11
rect 703 -19 704 -11
rect 706 -19 712 -11
rect 714 -19 715 -11
rect 733 -19 734 -11
rect 736 -19 742 -11
rect 744 -19 745 -11
rect 757 -19 758 -15
rect 760 -19 761 -15
rect 784 -19 785 -11
rect 787 -19 793 -11
rect 795 -19 796 -11
rect 808 -19 809 -15
rect 811 -19 812 -15
rect 830 -19 831 -11
rect 833 -19 834 -11
rect 838 -19 839 -11
rect 841 -19 842 -11
rect 854 -19 855 -15
rect 857 -19 858 -15
rect 889 -19 890 -15
rect 892 -19 893 -15
rect 907 -19 908 -15
rect 910 -19 911 -15
rect 925 -19 926 -11
rect 928 -19 934 -11
rect 936 -19 937 -11
rect 941 -19 942 -11
rect 944 -19 950 -11
rect 952 -19 953 -11
rect 970 -19 971 -15
rect 973 -19 974 -15
rect 988 -19 989 -15
rect 991 -19 992 -15
rect 1006 -19 1007 -11
rect 1009 -19 1015 -11
rect 1017 -19 1018 -11
rect 1022 -19 1023 -11
rect 1025 -19 1031 -11
rect 1033 -19 1034 -11
rect 1052 -19 1053 -11
rect 1055 -19 1061 -11
rect 1063 -19 1064 -11
rect 1076 -19 1077 -15
rect 1079 -19 1080 -15
rect 1103 -19 1104 -11
rect 1106 -19 1112 -11
rect 1114 -19 1115 -11
rect 1127 -19 1128 -15
rect 1130 -19 1131 -15
rect 1149 -19 1150 -11
rect 1152 -19 1153 -11
rect 1157 -19 1158 -11
rect 1160 -19 1161 -11
rect 1173 -19 1174 -15
rect 1176 -19 1177 -15
rect 1197 -19 1198 -15
rect 1200 -19 1201 -15
rect 1221 -19 1222 -15
rect 1224 -19 1225 -15
rect 1247 -19 1248 -15
rect 1250 -19 1251 -15
rect 1272 -19 1273 -15
rect 1275 -19 1276 -15
<< pdiffusion >>
rect -47 27 -46 35
rect -44 27 -43 35
rect -29 27 -28 35
rect -26 27 -25 35
rect -11 19 -10 35
rect -8 27 -7 35
rect -3 27 -2 35
rect -8 19 -2 27
rect 0 19 1 35
rect 5 19 6 35
rect 8 27 14 35
rect 8 19 9 27
rect 13 19 14 27
rect 16 19 17 35
rect 34 27 35 35
rect 37 27 38 35
rect 52 27 53 35
rect 55 27 56 35
rect 70 19 71 35
rect 73 27 74 35
rect 78 27 79 35
rect 73 19 79 27
rect 81 19 82 35
rect 86 19 87 35
rect 89 27 95 35
rect 89 19 90 27
rect 94 19 95 27
rect 97 19 98 35
rect 116 27 117 35
rect 119 27 120 35
rect 124 27 125 35
rect 127 27 128 35
rect 140 27 141 35
rect 143 27 144 35
rect 167 27 168 35
rect 170 27 171 35
rect 175 27 176 35
rect 178 27 179 35
rect 191 27 192 35
rect 194 27 195 35
rect 213 27 214 35
rect 216 27 222 35
rect 224 27 225 35
rect 237 27 238 35
rect 240 27 241 35
rect 261 27 262 35
rect 264 27 265 35
rect 279 27 280 35
rect 282 27 283 35
rect 297 19 298 35
rect 300 27 301 35
rect 305 27 306 35
rect 300 19 306 27
rect 308 19 309 35
rect 313 19 314 35
rect 316 27 322 35
rect 316 19 317 27
rect 321 19 322 27
rect 324 19 325 35
rect 342 27 343 35
rect 345 27 346 35
rect 360 27 361 35
rect 363 27 364 35
rect 378 19 379 35
rect 381 27 382 35
rect 386 27 387 35
rect 381 19 387 27
rect 389 19 390 35
rect 394 19 395 35
rect 397 27 403 35
rect 397 19 398 27
rect 402 19 403 27
rect 405 19 406 35
rect 424 27 425 35
rect 427 27 428 35
rect 432 27 433 35
rect 435 27 436 35
rect 448 27 449 35
rect 451 27 452 35
rect 475 27 476 35
rect 478 27 479 35
rect 483 27 484 35
rect 486 27 487 35
rect 499 27 500 35
rect 502 27 503 35
rect 521 27 522 35
rect 524 27 530 35
rect 532 27 533 35
rect 545 27 546 35
rect 548 27 549 35
rect 570 27 571 35
rect 573 27 574 35
rect 588 27 589 35
rect 591 27 592 35
rect 606 19 607 35
rect 609 27 610 35
rect 614 27 615 35
rect 609 19 615 27
rect 617 19 618 35
rect 622 19 623 35
rect 625 27 631 35
rect 625 19 626 27
rect 630 19 631 27
rect 633 19 634 35
rect 651 27 652 35
rect 654 27 655 35
rect 669 27 670 35
rect 672 27 673 35
rect 687 19 688 35
rect 690 27 691 35
rect 695 27 696 35
rect 690 19 696 27
rect 698 19 699 35
rect 703 19 704 35
rect 706 27 712 35
rect 706 19 707 27
rect 711 19 712 27
rect 714 19 715 35
rect 733 27 734 35
rect 736 27 737 35
rect 741 27 742 35
rect 744 27 745 35
rect 757 27 758 35
rect 760 27 761 35
rect 784 27 785 35
rect 787 27 788 35
rect 792 27 793 35
rect 795 27 796 35
rect 808 27 809 35
rect 811 27 812 35
rect 830 27 831 35
rect 833 27 839 35
rect 841 27 842 35
rect 854 27 855 35
rect 857 27 858 35
rect 889 27 890 35
rect 892 27 893 35
rect 907 27 908 35
rect 910 27 911 35
rect 925 19 926 35
rect 928 27 929 35
rect 933 27 934 35
rect 928 19 934 27
rect 936 19 937 35
rect 941 19 942 35
rect 944 27 950 35
rect 944 19 945 27
rect 949 19 950 27
rect 952 19 953 35
rect 970 27 971 35
rect 973 27 974 35
rect 988 27 989 35
rect 991 27 992 35
rect 1006 19 1007 35
rect 1009 27 1010 35
rect 1014 27 1015 35
rect 1009 19 1015 27
rect 1017 19 1018 35
rect 1022 19 1023 35
rect 1025 27 1031 35
rect 1025 19 1026 27
rect 1030 19 1031 27
rect 1033 19 1034 35
rect 1052 27 1053 35
rect 1055 27 1056 35
rect 1060 27 1061 35
rect 1063 27 1064 35
rect 1076 27 1077 35
rect 1079 27 1080 35
rect 1103 27 1104 35
rect 1106 27 1107 35
rect 1111 27 1112 35
rect 1114 27 1115 35
rect 1127 27 1128 35
rect 1130 27 1131 35
rect 1149 27 1150 35
rect 1152 27 1158 35
rect 1160 27 1161 35
rect 1173 27 1174 35
rect 1176 27 1177 35
rect 1197 27 1198 35
rect 1200 27 1201 35
rect 1221 27 1222 35
rect 1224 27 1225 35
rect 1247 27 1248 35
rect 1250 27 1251 35
rect 1272 27 1273 35
rect 1275 27 1276 35
<< metal1 >>
rect 56 84 175 88
rect 254 84 360 88
rect 364 84 483 88
rect 565 84 669 88
rect 673 84 792 88
rect 877 84 988 88
rect 992 84 1111 88
rect 38 77 167 81
rect 346 77 475 81
rect 655 77 784 81
rect 974 77 1103 81
rect -47 70 120 74
rect -47 51 -43 70
rect -29 58 -25 61
rect 116 59 120 70
rect 261 70 428 74
rect 124 59 128 62
rect -43 47 -11 51
rect 2 47 5 51
rect 41 47 70 51
rect 83 47 86 51
rect 261 51 265 70
rect 279 58 283 61
rect 424 59 428 70
rect 570 70 737 74
rect 432 59 436 62
rect 206 47 213 51
rect 265 47 297 51
rect 310 47 313 51
rect 349 47 378 51
rect 391 47 394 51
rect 570 51 574 70
rect 588 58 592 61
rect 733 59 737 70
rect 889 70 1056 74
rect 741 59 745 62
rect 514 47 521 51
rect 574 47 606 51
rect 619 47 622 51
rect 658 47 687 51
rect 700 47 703 51
rect 889 51 893 70
rect 907 58 911 61
rect 1052 59 1056 70
rect 1060 59 1064 62
rect 823 47 830 51
rect 893 47 925 51
rect 938 47 941 51
rect 977 47 1006 51
rect 1019 47 1022 51
rect 1142 47 1149 51
rect -51 43 1280 44
rect -51 39 -37 43
rect -33 39 46 43
rect 50 39 120 43
rect 124 39 137 43
rect 141 39 171 43
rect 175 39 188 43
rect 192 39 217 43
rect 221 39 234 43
rect 238 39 271 43
rect 275 39 354 43
rect 358 39 428 43
rect 432 39 445 43
rect 449 39 479 43
rect 483 39 496 43
rect 500 39 525 43
rect 529 39 542 43
rect 546 39 580 43
rect 584 39 663 43
rect 667 39 737 43
rect 741 39 754 43
rect 758 39 788 43
rect 792 39 805 43
rect 809 39 834 43
rect 838 39 851 43
rect 855 39 899 43
rect 903 39 982 43
rect 986 39 1056 43
rect 1060 39 1073 43
rect 1077 39 1107 43
rect 1111 39 1124 43
rect 1128 39 1153 43
rect 1157 39 1170 43
rect 1174 39 1194 43
rect 1198 39 1218 43
rect 1222 39 1244 43
rect 1248 39 1269 43
rect 1273 39 1280 43
rect -51 38 1280 39
rect -51 35 -47 38
rect -33 35 -29 38
rect -7 35 -3 38
rect 30 35 34 38
rect 48 35 52 38
rect 74 35 78 38
rect 112 35 116 38
rect 128 35 132 38
rect -43 12 -39 27
rect -25 12 -21 27
rect -11 19 1 23
rect 5 31 17 35
rect 9 7 13 19
rect 38 12 42 27
rect 56 12 60 27
rect 70 19 82 23
rect 86 31 98 35
rect 136 35 140 38
rect 163 35 167 38
rect 179 35 183 38
rect 187 35 191 38
rect 209 35 213 38
rect 233 35 237 38
rect 257 35 261 38
rect 275 35 279 38
rect 301 35 305 38
rect 338 35 342 38
rect 356 35 360 38
rect 382 35 386 38
rect 420 35 424 38
rect 436 35 440 38
rect 90 7 94 19
rect 120 12 124 27
rect 144 12 148 27
rect 171 12 175 27
rect 195 12 199 27
rect 225 12 229 27
rect 241 12 245 27
rect 265 12 269 27
rect 283 12 287 27
rect 297 19 309 23
rect 313 31 325 35
rect 120 8 137 12
rect -43 -15 -39 7
rect -25 -15 -21 7
rect 1 3 31 7
rect 1 -11 5 3
rect 38 -15 42 7
rect 56 -15 60 7
rect 82 3 104 7
rect 82 -11 86 3
rect 128 -11 132 8
rect -51 -22 -47 -19
rect -33 -22 -29 -19
rect -15 -22 -11 -19
rect 17 -22 21 -19
rect 30 -22 34 -19
rect 48 -22 52 -19
rect 66 -22 70 -19
rect 98 -22 102 -19
rect 171 8 188 12
rect 144 -15 148 7
rect 179 -11 183 8
rect 217 8 234 12
rect 241 8 249 12
rect 195 -15 199 7
rect 217 -11 221 8
rect 241 -15 245 8
rect 317 7 321 19
rect 346 12 350 27
rect 364 12 368 27
rect 378 19 390 23
rect 394 31 406 35
rect 444 35 448 38
rect 471 35 475 38
rect 487 35 491 38
rect 495 35 499 38
rect 517 35 521 38
rect 541 35 545 38
rect 566 35 570 38
rect 584 35 588 38
rect 610 35 614 38
rect 647 35 651 38
rect 665 35 669 38
rect 691 35 695 38
rect 729 35 733 38
rect 745 35 749 38
rect 398 7 402 19
rect 428 12 432 27
rect 452 12 456 27
rect 479 12 483 27
rect 503 12 507 27
rect 533 12 537 27
rect 549 12 553 27
rect 428 8 445 12
rect 265 -15 269 7
rect 283 -15 287 7
rect 309 3 339 7
rect 309 -11 313 3
rect 112 -22 116 -19
rect 136 -22 140 -19
rect 163 -22 167 -19
rect 187 -22 191 -19
rect 209 -22 213 -19
rect 225 -22 229 -19
rect 346 -15 350 7
rect 364 -15 368 7
rect 390 3 412 7
rect 390 -11 394 3
rect 436 -11 440 8
rect 233 -22 237 -19
rect 257 -22 261 -19
rect 275 -22 279 -19
rect 293 -22 297 -19
rect 325 -22 329 -19
rect 338 -22 342 -19
rect 356 -22 360 -19
rect 374 -22 378 -19
rect 406 -22 410 -19
rect 479 8 496 12
rect 452 -15 456 7
rect 487 -11 491 8
rect 525 8 542 12
rect 549 8 559 12
rect 574 12 578 27
rect 592 12 596 27
rect 606 19 618 23
rect 622 31 634 35
rect 503 -15 507 7
rect 525 -11 529 8
rect 549 -15 553 8
rect 626 7 630 19
rect 655 12 659 27
rect 673 12 677 27
rect 687 19 699 23
rect 703 31 715 35
rect 753 35 757 38
rect 780 35 784 38
rect 796 35 800 38
rect 804 35 808 38
rect 826 35 830 38
rect 850 35 854 38
rect 885 35 889 38
rect 903 35 907 38
rect 929 35 933 38
rect 966 35 970 38
rect 984 35 988 38
rect 1010 35 1014 38
rect 1048 35 1052 38
rect 1064 35 1068 38
rect 707 7 711 19
rect 737 12 741 27
rect 761 12 765 27
rect 788 12 792 27
rect 812 12 816 27
rect 842 12 846 27
rect 858 12 862 27
rect 737 8 754 12
rect 574 -15 578 7
rect 592 -15 596 7
rect 618 3 648 7
rect 618 -11 622 3
rect 420 -22 424 -19
rect 444 -22 448 -19
rect 471 -22 475 -19
rect 495 -22 499 -19
rect 517 -22 521 -19
rect 533 -22 537 -19
rect 655 -15 659 7
rect 673 -15 677 7
rect 699 3 721 7
rect 699 -11 703 3
rect 745 -11 749 8
rect 541 -22 545 -19
rect 566 -22 570 -19
rect 584 -22 588 -19
rect 602 -22 606 -19
rect 634 -22 638 -19
rect 647 -22 651 -19
rect 665 -22 669 -19
rect 683 -22 687 -19
rect 715 -22 719 -19
rect 788 8 805 12
rect 761 -15 765 7
rect 796 -11 800 8
rect 834 8 851 12
rect 858 8 872 12
rect 893 12 897 27
rect 911 12 915 27
rect 925 19 937 23
rect 941 31 953 35
rect 812 -15 816 7
rect 834 -11 838 8
rect 858 -15 862 8
rect 945 7 949 19
rect 974 12 978 27
rect 992 12 996 27
rect 1006 19 1018 23
rect 1022 31 1034 35
rect 1072 35 1076 38
rect 1099 35 1103 38
rect 1115 35 1119 38
rect 1123 35 1127 38
rect 1145 35 1149 38
rect 1169 35 1173 38
rect 1193 35 1197 38
rect 1217 35 1221 38
rect 1243 35 1247 38
rect 1268 35 1272 38
rect 1026 7 1030 19
rect 1056 12 1060 27
rect 1080 12 1084 27
rect 1107 12 1111 27
rect 1131 12 1135 27
rect 1161 12 1165 27
rect 1177 12 1181 27
rect 1201 12 1205 27
rect 1056 8 1073 12
rect 893 -15 897 7
rect 911 -15 915 7
rect 937 3 967 7
rect 937 -11 941 3
rect 729 -22 733 -19
rect 753 -22 757 -19
rect 780 -22 784 -19
rect 804 -22 808 -19
rect 826 -22 830 -19
rect 842 -22 846 -19
rect 974 -15 978 7
rect 992 -15 996 7
rect 1018 3 1040 7
rect 1018 -11 1022 3
rect 1064 -11 1068 8
rect 850 -22 854 -19
rect 885 -22 889 -19
rect 903 -22 907 -19
rect 921 -22 925 -19
rect 953 -22 957 -19
rect 966 -22 970 -19
rect 984 -22 988 -19
rect 1002 -22 1006 -19
rect 1034 -22 1038 -19
rect 1107 8 1124 12
rect 1080 -15 1084 7
rect 1115 -11 1119 8
rect 1153 8 1170 12
rect 1177 8 1194 12
rect 1201 8 1218 12
rect 1131 -15 1135 7
rect 1153 -11 1157 8
rect 1177 -15 1181 8
rect 1201 -15 1205 8
rect 1225 -15 1229 27
rect 1251 12 1255 27
rect 1048 -22 1052 -19
rect 1072 -22 1076 -19
rect 1099 -22 1103 -19
rect 1123 -22 1127 -19
rect 1145 -22 1149 -19
rect 1161 -22 1165 -19
rect 1236 8 1244 12
rect 1251 8 1269 12
rect 1169 -22 1173 -19
rect 1193 -22 1197 -19
rect 1217 -22 1221 -19
rect -51 -23 1227 -22
rect -51 -27 -50 -23
rect -46 -27 31 -23
rect 35 -27 113 -23
rect 117 -27 137 -23
rect 141 -27 164 -23
rect 168 -27 188 -23
rect 192 -27 210 -23
rect 214 -27 234 -23
rect 238 -27 258 -23
rect 262 -27 339 -23
rect 343 -27 421 -23
rect 425 -27 445 -23
rect 449 -27 472 -23
rect 476 -27 496 -23
rect 500 -27 518 -23
rect 522 -27 542 -23
rect 546 -27 567 -23
rect 571 -27 648 -23
rect 652 -27 730 -23
rect 734 -27 754 -23
rect 758 -27 781 -23
rect 785 -27 805 -23
rect 809 -27 827 -23
rect 831 -27 851 -23
rect 855 -27 886 -23
rect 890 -27 967 -23
rect 971 -27 1049 -23
rect 1053 -27 1073 -23
rect 1077 -27 1100 -23
rect 1104 -27 1124 -23
rect 1128 -27 1146 -23
rect 1150 -27 1170 -23
rect 1174 -27 1194 -23
rect 1198 -27 1218 -23
rect 1222 -27 1227 -23
rect -51 -28 1227 -27
rect -25 -35 -3 -31
rect 10 -35 13 -31
rect 56 -35 78 -31
rect 91 -35 94 -31
rect 217 -35 221 -31
rect 283 -35 305 -31
rect 318 -35 321 -31
rect 364 -35 386 -31
rect 399 -35 402 -31
rect 525 -35 529 -31
rect 592 -35 614 -31
rect 627 -35 630 -31
rect 673 -35 695 -31
rect 708 -35 711 -31
rect 834 -35 838 -31
rect 911 -35 933 -31
rect 946 -35 949 -31
rect 992 -35 1014 -31
rect 1027 -35 1030 -31
rect 1153 -35 1157 -31
rect 1236 -52 1240 8
rect 1251 -15 1255 8
rect 1276 -15 1280 27
rect 1243 -22 1247 -19
rect 1268 -22 1272 -19
rect 1243 -23 1258 -22
rect 1243 -27 1244 -23
rect 1248 -27 1258 -23
rect 1243 -28 1258 -27
rect 1264 -23 1280 -22
rect 1264 -27 1269 -23
rect 1273 -27 1280 -23
rect 1264 -28 1280 -27
rect 1044 -56 1240 -52
<< metal2 >>
rect -24 62 124 66
rect -3 44 1 47
rect 78 44 82 47
rect 201 44 205 47
rect -24 40 1 44
rect 57 40 82 44
rect 145 40 205 44
rect -24 12 -20 40
rect 57 12 61 40
rect 145 12 149 40
rect 250 12 254 84
rect 284 62 432 66
rect 305 44 309 47
rect 386 44 390 47
rect 509 44 513 47
rect 284 40 309 44
rect 365 40 390 44
rect 453 40 513 44
rect 284 12 288 40
rect 365 12 369 40
rect 453 12 457 40
rect 560 13 564 84
rect 593 62 741 66
rect 614 44 618 47
rect 695 44 699 47
rect 818 44 822 47
rect 593 40 618 44
rect 674 40 699 44
rect 762 40 822 44
rect 593 12 597 40
rect 674 12 678 40
rect 762 12 766 40
rect 873 13 877 84
rect 912 62 1060 66
rect 933 44 937 47
rect 1014 44 1018 47
rect 1137 44 1141 47
rect 912 40 937 44
rect 993 40 1018 44
rect 1081 40 1141 44
rect 912 12 916 40
rect 993 12 997 40
rect 1081 12 1085 40
rect -42 -24 -38 7
rect 39 -24 43 7
rect -42 -28 9 -24
rect 39 -28 90 -24
rect 5 -31 9 -28
rect 86 -31 90 -28
rect 196 -31 200 7
rect 266 -24 270 7
rect 347 -24 351 7
rect 266 -28 317 -24
rect 347 -28 398 -24
rect 313 -31 317 -28
rect 394 -31 398 -28
rect 504 -31 508 7
rect 575 -24 579 7
rect 656 -24 660 7
rect 575 -28 626 -24
rect 656 -28 707 -24
rect 622 -31 626 -28
rect 703 -31 707 -28
rect 813 -31 817 7
rect 894 -24 898 7
rect 975 -24 979 7
rect 894 -28 945 -24
rect 975 -28 1026 -24
rect 941 -31 945 -28
rect 1022 -31 1026 -28
rect 196 -35 212 -31
rect 504 -35 520 -31
rect 813 -35 829 -31
rect 1040 -52 1044 3
rect 1132 -31 1136 7
rect 1132 -35 1148 -31
rect 1227 -34 1233 -28
rect 1258 -34 1264 -28
rect 1227 -40 1264 -34
<< ntransistor >>
rect -46 -19 -44 -15
rect -28 -19 -26 -15
rect -10 -19 -8 -11
rect -2 -19 0 -11
rect 6 -19 8 -11
rect 14 -19 16 -11
rect 35 -19 37 -15
rect 53 -19 55 -15
rect 71 -19 73 -11
rect 79 -19 81 -11
rect 87 -19 89 -11
rect 95 -19 97 -11
rect 117 -19 119 -11
rect 125 -19 127 -11
rect 141 -19 143 -15
rect 168 -19 170 -11
rect 176 -19 178 -11
rect 192 -19 194 -15
rect 214 -19 216 -11
rect 222 -19 224 -11
rect 238 -19 240 -15
rect 262 -19 264 -15
rect 280 -19 282 -15
rect 298 -19 300 -11
rect 306 -19 308 -11
rect 314 -19 316 -11
rect 322 -19 324 -11
rect 343 -19 345 -15
rect 361 -19 363 -15
rect 379 -19 381 -11
rect 387 -19 389 -11
rect 395 -19 397 -11
rect 403 -19 405 -11
rect 425 -19 427 -11
rect 433 -19 435 -11
rect 449 -19 451 -15
rect 476 -19 478 -11
rect 484 -19 486 -11
rect 500 -19 502 -15
rect 522 -19 524 -11
rect 530 -19 532 -11
rect 546 -19 548 -15
rect 571 -19 573 -15
rect 589 -19 591 -15
rect 607 -19 609 -11
rect 615 -19 617 -11
rect 623 -19 625 -11
rect 631 -19 633 -11
rect 652 -19 654 -15
rect 670 -19 672 -15
rect 688 -19 690 -11
rect 696 -19 698 -11
rect 704 -19 706 -11
rect 712 -19 714 -11
rect 734 -19 736 -11
rect 742 -19 744 -11
rect 758 -19 760 -15
rect 785 -19 787 -11
rect 793 -19 795 -11
rect 809 -19 811 -15
rect 831 -19 833 -11
rect 839 -19 841 -11
rect 855 -19 857 -15
rect 890 -19 892 -15
rect 908 -19 910 -15
rect 926 -19 928 -11
rect 934 -19 936 -11
rect 942 -19 944 -11
rect 950 -19 952 -11
rect 971 -19 973 -15
rect 989 -19 991 -15
rect 1007 -19 1009 -11
rect 1015 -19 1017 -11
rect 1023 -19 1025 -11
rect 1031 -19 1033 -11
rect 1053 -19 1055 -11
rect 1061 -19 1063 -11
rect 1077 -19 1079 -15
rect 1104 -19 1106 -11
rect 1112 -19 1114 -11
rect 1128 -19 1130 -15
rect 1150 -19 1152 -11
rect 1158 -19 1160 -11
rect 1174 -19 1176 -15
rect 1198 -19 1200 -15
rect 1222 -19 1224 -15
rect 1248 -19 1250 -15
rect 1273 -19 1275 -15
<< ptransistor >>
rect -46 27 -44 35
rect -28 27 -26 35
rect -10 19 -8 35
rect -2 19 0 35
rect 6 19 8 35
rect 14 19 16 35
rect 35 27 37 35
rect 53 27 55 35
rect 71 19 73 35
rect 79 19 81 35
rect 87 19 89 35
rect 95 19 97 35
rect 117 27 119 35
rect 125 27 127 35
rect 141 27 143 35
rect 168 27 170 35
rect 176 27 178 35
rect 192 27 194 35
rect 214 27 216 35
rect 222 27 224 35
rect 238 27 240 35
rect 262 27 264 35
rect 280 27 282 35
rect 298 19 300 35
rect 306 19 308 35
rect 314 19 316 35
rect 322 19 324 35
rect 343 27 345 35
rect 361 27 363 35
rect 379 19 381 35
rect 387 19 389 35
rect 395 19 397 35
rect 403 19 405 35
rect 425 27 427 35
rect 433 27 435 35
rect 449 27 451 35
rect 476 27 478 35
rect 484 27 486 35
rect 500 27 502 35
rect 522 27 524 35
rect 530 27 532 35
rect 546 27 548 35
rect 571 27 573 35
rect 589 27 591 35
rect 607 19 609 35
rect 615 19 617 35
rect 623 19 625 35
rect 631 19 633 35
rect 652 27 654 35
rect 670 27 672 35
rect 688 19 690 35
rect 696 19 698 35
rect 704 19 706 35
rect 712 19 714 35
rect 734 27 736 35
rect 742 27 744 35
rect 758 27 760 35
rect 785 27 787 35
rect 793 27 795 35
rect 809 27 811 35
rect 831 27 833 35
rect 839 27 841 35
rect 855 27 857 35
rect 890 27 892 35
rect 908 27 910 35
rect 926 19 928 35
rect 934 19 936 35
rect 942 19 944 35
rect 950 19 952 35
rect 971 27 973 35
rect 989 27 991 35
rect 1007 19 1009 35
rect 1015 19 1017 35
rect 1023 19 1025 35
rect 1031 19 1033 35
rect 1053 27 1055 35
rect 1061 27 1063 35
rect 1077 27 1079 35
rect 1104 27 1106 35
rect 1112 27 1114 35
rect 1128 27 1130 35
rect 1150 27 1152 35
rect 1158 27 1160 35
rect 1174 27 1176 35
rect 1198 27 1200 35
rect 1222 27 1224 35
rect 1248 27 1250 35
rect 1273 27 1275 35
<< polycontact >>
rect 52 84 56 88
rect 175 84 179 88
rect 360 84 364 88
rect 483 84 487 88
rect 669 84 673 88
rect 792 84 796 88
rect 988 84 992 88
rect 1111 84 1115 88
rect 34 77 38 81
rect -29 54 -25 58
rect -47 47 -43 51
rect -11 47 -7 51
rect 5 47 9 51
rect 37 47 41 51
rect 167 77 171 81
rect 116 55 120 59
rect 124 55 128 59
rect 70 47 74 51
rect 86 47 90 51
rect 342 77 346 81
rect 279 54 283 58
rect 213 47 217 51
rect 261 47 265 51
rect 297 47 301 51
rect 313 47 317 51
rect 345 47 349 51
rect 475 77 479 81
rect 424 55 428 59
rect 432 55 436 59
rect 378 47 382 51
rect 394 47 398 51
rect 651 77 655 81
rect 588 54 592 58
rect 521 47 525 51
rect 570 47 574 51
rect 606 47 610 51
rect 622 47 626 51
rect 654 47 658 51
rect 784 77 788 81
rect 733 55 737 59
rect 741 55 745 59
rect 687 47 691 51
rect 703 47 707 51
rect 970 77 974 81
rect 907 54 911 58
rect 830 47 834 51
rect 889 47 893 51
rect 925 47 929 51
rect 941 47 945 51
rect 973 47 977 51
rect 1103 77 1107 81
rect 1052 55 1056 59
rect 1060 55 1064 59
rect 1006 47 1010 51
rect 1022 47 1026 51
rect 1149 47 1153 51
rect -32 8 -28 12
rect 31 3 35 7
rect 137 8 141 12
rect 188 8 192 12
rect 234 8 238 12
rect 276 8 280 12
rect 339 3 343 7
rect 445 8 449 12
rect 496 8 500 12
rect 542 8 546 12
rect 585 8 589 12
rect 648 3 652 7
rect 754 8 758 12
rect 805 8 809 12
rect 851 8 855 12
rect 904 8 908 12
rect 967 3 971 7
rect 1073 8 1077 12
rect 1124 8 1128 12
rect 1170 8 1174 12
rect 1194 8 1198 12
rect 1218 8 1222 12
rect 1244 8 1248 12
rect 1269 8 1273 12
rect -29 -35 -25 -31
rect -3 -35 1 -31
rect 13 -35 17 -31
rect 52 -35 56 -31
rect 78 -35 82 -31
rect 94 -35 98 -31
rect 221 -35 225 -31
rect 279 -35 283 -31
rect 305 -35 309 -31
rect 321 -35 325 -31
rect 360 -35 364 -31
rect 386 -35 390 -31
rect 402 -35 406 -31
rect 529 -35 533 -31
rect 588 -35 592 -31
rect 614 -35 618 -31
rect 630 -35 634 -31
rect 669 -35 673 -31
rect 695 -35 699 -31
rect 711 -35 715 -31
rect 838 -35 842 -31
rect 907 -35 911 -31
rect 933 -35 937 -31
rect 949 -35 953 -31
rect 988 -35 992 -31
rect 1014 -35 1018 -31
rect 1030 -35 1034 -31
rect 1157 -35 1161 -31
<< ndcontact >>
rect -51 -19 -47 -15
rect -43 -19 -39 -15
rect -33 -19 -29 -15
rect -25 -19 -21 -15
rect -15 -19 -11 -11
rect 1 -19 5 -11
rect 17 -19 21 -11
rect 30 -19 34 -15
rect 38 -19 42 -15
rect 48 -19 52 -15
rect 56 -19 60 -15
rect 66 -19 70 -11
rect 82 -19 86 -11
rect 98 -19 102 -11
rect 112 -19 116 -11
rect 128 -19 132 -11
rect 136 -19 140 -15
rect 144 -19 148 -15
rect 163 -19 167 -11
rect 179 -19 183 -11
rect 187 -19 191 -15
rect 195 -19 199 -15
rect 209 -19 213 -11
rect 217 -19 221 -11
rect 225 -19 229 -11
rect 233 -19 237 -15
rect 241 -19 245 -15
rect 257 -19 261 -15
rect 265 -19 269 -15
rect 275 -19 279 -15
rect 283 -19 287 -15
rect 293 -19 297 -11
rect 309 -19 313 -11
rect 325 -19 329 -11
rect 338 -19 342 -15
rect 346 -19 350 -15
rect 356 -19 360 -15
rect 364 -19 368 -15
rect 374 -19 378 -11
rect 390 -19 394 -11
rect 406 -19 410 -11
rect 420 -19 424 -11
rect 436 -19 440 -11
rect 444 -19 448 -15
rect 452 -19 456 -15
rect 471 -19 475 -11
rect 487 -19 491 -11
rect 495 -19 499 -15
rect 503 -19 507 -15
rect 517 -19 521 -11
rect 525 -19 529 -11
rect 533 -19 537 -11
rect 541 -19 545 -15
rect 549 -19 553 -15
rect 566 -19 570 -15
rect 574 -19 578 -15
rect 584 -19 588 -15
rect 592 -19 596 -15
rect 602 -19 606 -11
rect 618 -19 622 -11
rect 634 -19 638 -11
rect 647 -19 651 -15
rect 655 -19 659 -15
rect 665 -19 669 -15
rect 673 -19 677 -15
rect 683 -19 687 -11
rect 699 -19 703 -11
rect 715 -19 719 -11
rect 729 -19 733 -11
rect 745 -19 749 -11
rect 753 -19 757 -15
rect 761 -19 765 -15
rect 780 -19 784 -11
rect 796 -19 800 -11
rect 804 -19 808 -15
rect 812 -19 816 -15
rect 826 -19 830 -11
rect 834 -19 838 -11
rect 842 -19 846 -11
rect 850 -19 854 -15
rect 858 -19 862 -15
rect 885 -19 889 -15
rect 893 -19 897 -15
rect 903 -19 907 -15
rect 911 -19 915 -15
rect 921 -19 925 -11
rect 937 -19 941 -11
rect 953 -19 957 -11
rect 966 -19 970 -15
rect 974 -19 978 -15
rect 984 -19 988 -15
rect 992 -19 996 -15
rect 1002 -19 1006 -11
rect 1018 -19 1022 -11
rect 1034 -19 1038 -11
rect 1048 -19 1052 -11
rect 1064 -19 1068 -11
rect 1072 -19 1076 -15
rect 1080 -19 1084 -15
rect 1099 -19 1103 -11
rect 1115 -19 1119 -11
rect 1123 -19 1127 -15
rect 1131 -19 1135 -15
rect 1145 -19 1149 -11
rect 1153 -19 1157 -11
rect 1161 -19 1165 -11
rect 1169 -19 1173 -15
rect 1177 -19 1181 -15
rect 1193 -19 1197 -15
rect 1201 -19 1205 -15
rect 1217 -19 1221 -15
rect 1225 -19 1229 -15
rect 1243 -19 1247 -15
rect 1251 -19 1255 -15
rect 1268 -19 1272 -15
rect 1276 -19 1280 -15
<< pdcontact >>
rect -51 27 -47 35
rect -43 27 -39 35
rect -33 27 -29 35
rect -25 27 -21 35
rect -15 19 -11 35
rect -7 27 -3 35
rect 1 19 5 35
rect 9 19 13 27
rect 17 19 21 35
rect 30 27 34 35
rect 38 27 42 35
rect 48 27 52 35
rect 56 27 60 35
rect 66 19 70 35
rect 74 27 78 35
rect 82 19 86 35
rect 90 19 94 27
rect 98 19 102 35
rect 112 27 116 35
rect 120 27 124 35
rect 128 27 132 35
rect 136 27 140 35
rect 144 27 148 35
rect 163 27 167 35
rect 171 27 175 35
rect 179 27 183 35
rect 187 27 191 35
rect 195 27 199 35
rect 209 27 213 35
rect 225 27 229 35
rect 233 27 237 35
rect 241 27 245 35
rect 257 27 261 35
rect 265 27 269 35
rect 275 27 279 35
rect 283 27 287 35
rect 293 19 297 35
rect 301 27 305 35
rect 309 19 313 35
rect 317 19 321 27
rect 325 19 329 35
rect 338 27 342 35
rect 346 27 350 35
rect 356 27 360 35
rect 364 27 368 35
rect 374 19 378 35
rect 382 27 386 35
rect 390 19 394 35
rect 398 19 402 27
rect 406 19 410 35
rect 420 27 424 35
rect 428 27 432 35
rect 436 27 440 35
rect 444 27 448 35
rect 452 27 456 35
rect 471 27 475 35
rect 479 27 483 35
rect 487 27 491 35
rect 495 27 499 35
rect 503 27 507 35
rect 517 27 521 35
rect 533 27 537 35
rect 541 27 545 35
rect 549 27 553 35
rect 566 27 570 35
rect 574 27 578 35
rect 584 27 588 35
rect 592 27 596 35
rect 602 19 606 35
rect 610 27 614 35
rect 618 19 622 35
rect 626 19 630 27
rect 634 19 638 35
rect 647 27 651 35
rect 655 27 659 35
rect 665 27 669 35
rect 673 27 677 35
rect 683 19 687 35
rect 691 27 695 35
rect 699 19 703 35
rect 707 19 711 27
rect 715 19 719 35
rect 729 27 733 35
rect 737 27 741 35
rect 745 27 749 35
rect 753 27 757 35
rect 761 27 765 35
rect 780 27 784 35
rect 788 27 792 35
rect 796 27 800 35
rect 804 27 808 35
rect 812 27 816 35
rect 826 27 830 35
rect 842 27 846 35
rect 850 27 854 35
rect 858 27 862 35
rect 885 27 889 35
rect 893 27 897 35
rect 903 27 907 35
rect 911 27 915 35
rect 921 19 925 35
rect 929 27 933 35
rect 937 19 941 35
rect 945 19 949 27
rect 953 19 957 35
rect 966 27 970 35
rect 974 27 978 35
rect 984 27 988 35
rect 992 27 996 35
rect 1002 19 1006 35
rect 1010 27 1014 35
rect 1018 19 1022 35
rect 1026 19 1030 27
rect 1034 19 1038 35
rect 1048 27 1052 35
rect 1056 27 1060 35
rect 1064 27 1068 35
rect 1072 27 1076 35
rect 1080 27 1084 35
rect 1099 27 1103 35
rect 1107 27 1111 35
rect 1115 27 1119 35
rect 1123 27 1127 35
rect 1131 27 1135 35
rect 1145 27 1149 35
rect 1161 27 1165 35
rect 1169 27 1173 35
rect 1177 27 1181 35
rect 1193 27 1197 35
rect 1201 27 1205 35
rect 1217 27 1221 35
rect 1225 27 1229 35
rect 1243 27 1247 35
rect 1251 27 1255 35
rect 1268 27 1272 35
rect 1276 27 1280 35
<< m2contact >>
rect 249 84 254 89
rect 560 84 565 89
rect 872 84 877 89
rect -29 61 -24 66
rect 124 62 129 67
rect -3 47 2 52
rect 78 47 83 52
rect 201 47 206 52
rect 279 61 284 66
rect 432 62 437 67
rect 305 47 310 52
rect 386 47 391 52
rect 509 47 514 52
rect 588 61 593 66
rect 741 62 746 67
rect 614 47 619 52
rect 695 47 700 52
rect 818 47 823 52
rect 907 61 912 66
rect 1060 62 1065 67
rect 933 47 938 52
rect 1014 47 1019 52
rect 1137 47 1142 52
rect -43 7 -38 12
rect -25 7 -20 12
rect 38 7 43 12
rect 56 7 61 12
rect 144 7 149 12
rect 195 7 200 12
rect 249 7 254 12
rect 265 7 270 12
rect 283 7 288 12
rect 346 7 351 12
rect 364 7 369 12
rect 452 7 457 12
rect 503 7 508 12
rect 559 8 564 13
rect 574 7 579 12
rect 592 7 597 12
rect 655 7 660 12
rect 673 7 678 12
rect 761 7 766 12
rect 812 7 817 12
rect 872 8 877 13
rect 893 7 898 12
rect 911 7 916 12
rect 974 7 979 12
rect 992 7 997 12
rect 1040 3 1044 7
rect 1080 7 1085 12
rect 1131 7 1136 12
rect 1227 -28 1233 -22
rect 5 -36 10 -31
rect 86 -36 91 -31
rect 212 -36 217 -31
rect 313 -36 318 -31
rect 394 -36 399 -31
rect 520 -36 525 -31
rect 622 -36 627 -31
rect 703 -36 708 -31
rect 829 -36 834 -31
rect 941 -36 946 -31
rect 1022 -36 1027 -31
rect 1148 -36 1153 -31
rect 1258 -28 1264 -22
rect 1040 -56 1044 -52
<< psubstratepcontact >>
rect -50 -27 -46 -23
rect 31 -27 35 -23
rect 113 -27 117 -23
rect 137 -27 141 -23
rect 164 -27 168 -23
rect 188 -27 192 -23
rect 210 -27 214 -23
rect 234 -27 238 -23
rect 258 -27 262 -23
rect 339 -27 343 -23
rect 421 -27 425 -23
rect 445 -27 449 -23
rect 472 -27 476 -23
rect 496 -27 500 -23
rect 518 -27 522 -23
rect 542 -27 546 -23
rect 567 -27 571 -23
rect 648 -27 652 -23
rect 730 -27 734 -23
rect 754 -27 758 -23
rect 781 -27 785 -23
rect 805 -27 809 -23
rect 827 -27 831 -23
rect 851 -27 855 -23
rect 886 -27 890 -23
rect 967 -27 971 -23
rect 1049 -27 1053 -23
rect 1073 -27 1077 -23
rect 1100 -27 1104 -23
rect 1124 -27 1128 -23
rect 1146 -27 1150 -23
rect 1170 -27 1174 -23
rect 1194 -27 1198 -23
rect 1218 -27 1222 -23
rect 1244 -27 1248 -23
rect 1269 -27 1273 -23
<< nsubstratencontact >>
rect -37 39 -33 43
rect 46 39 50 43
rect 120 39 124 43
rect 137 39 141 43
rect 171 39 175 43
rect 188 39 192 43
rect 217 39 221 43
rect 234 39 238 43
rect 271 39 275 43
rect 354 39 358 43
rect 428 39 432 43
rect 445 39 449 43
rect 479 39 483 43
rect 496 39 500 43
rect 525 39 529 43
rect 542 39 546 43
rect 580 39 584 43
rect 663 39 667 43
rect 737 39 741 43
rect 754 39 758 43
rect 788 39 792 43
rect 805 39 809 43
rect 834 39 838 43
rect 851 39 855 43
rect 899 39 903 43
rect 982 39 986 43
rect 1056 39 1060 43
rect 1073 39 1077 43
rect 1107 39 1111 43
rect 1124 39 1128 43
rect 1153 39 1157 43
rect 1170 39 1174 43
rect 1194 39 1198 43
rect 1218 39 1222 43
rect 1244 39 1248 43
rect 1269 39 1273 43
<< labels >>
rlabel polycontact -45 49 -45 49 1 A1
rlabel polycontact -30 10 -30 10 1 B1
rlabel metal1 25 41 25 41 1 vdd
rlabel metal1 25 -24 25 -24 1 gnd
rlabel polycontact 54 86 54 86 5 cin
rlabel metal1 101 5 101 5 1 S1
rlabel metal1 245 10 245 10 1 cout1
rlabel polycontact 263 49 263 49 1 A2
rlabel polycontact 278 10 278 10 1 B2
rlabel polycontact 362 86 362 86 5 cin2
rlabel metal1 409 5 409 5 1 S2
rlabel metal1 551 10 551 10 7 cout2
rlabel polycontact 572 49 572 49 1 A3
rlabel polycontact 587 10 587 10 1 B3
rlabel polycontact 671 86 671 86 5 cin3
rlabel metal1 719 5 719 5 1 S3
rlabel metal1 860 10 860 10 7 cout3
rlabel polycontact 891 49 891 49 1 A4
rlabel polycontact 906 10 906 10 1 B4
rlabel polycontact 990 86 990 86 5 cin4
rlabel metal1 1037 5 1037 5 1 S4
rlabel metal1 1179 10 1179 10 7 cout4
rlabel metal1 1227 10 1227 10 7 cout
rlabel metal1 1278 10 1278 10 7 sum
<< end >>
